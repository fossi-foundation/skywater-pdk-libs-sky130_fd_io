* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Placeholder for "condiode", which probably represents the parasitic
* well-to-substrate diode, although it does not take any parameters.
.SUBCKT sky130_fd_io__condiode NEG POS
.ENDS

.SUBCKT sky130_fd_io__gnd2gnd_120x2_lv_isosub BDY2_B2B SRC_BDY_LVC1 VSSD
XD0 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 area=90E+12 perim=132E+6
XD1 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 area=90E+12 perim=132E+6
.ENDS

.SUBCKT sky130_fd_io__amuxsplitv2_delay ENABLE_VDDA_H HLD_VDDA_H_N HOLD RESET
+ VCC_IO VGND
*.PININFO ENABLE_VDDA_H:I HLD_VDDA_H_N:I HOLD:O RESET:O VCC_IO:B
*.PININFO VGND:B
XI33 enable_vdda_switch hld_vdda_h_n_switch RESET VGND VCC_IO
+ sky130_fd_io__hvsbt_nand2
XI29 hld_vdda_h_n_switch hld_vdda_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI28 hld_vdda_h HLD_VDDA_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI12 enable_vdda_switch enable_vdda_h_n VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI13 enable_vdda_h_n ENABLE_VDDA_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI36 HOLD RESET VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 hld_vdda_h_n_switch hld_vdda_h VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2
+ w=1.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI30 hld_vdda_h HLD_VDDA_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 enable_vdda_switch enable_vdda_h_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5
+ m=2 w=1.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI15 enable_vdda_h_n ENABLE_VDDA_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI37 HOLD RESET VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_delay

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch AMUXBUS_L AMUXBUS_R NGATE_SL_H
+ NGATE_SR_H NMID_H PGATE_SL_H_N PGATE_SR_H_N VDDA VSSA
*.PININFO AMUXBUS_L:B AMUXBUS_R:B NGATE_SL_H:I NGATE_SR_H:I NMID_H:I
*.PININFO PGATE_SL_H_N:I PGATE_SR_H_N:I VDDA:B VSSA:B
xI20 mid VDDA sky130_fd_io__condiode
xI19 VSSA VDDA sky130_fd_io__condiode
XI18 VSSA nmid_h_s sky130_fd_io__res75only_small
XI1 AMUXBUS_L NGATE_SL_H mid mid sky130_fd_pr__nfet_g5v0d10v5 m=30 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 mid NGATE_SR_H AMUXBUS_R mid sky130_fd_pr__nfet_g5v0d10v5 m=30 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 mid NMID_H nmid_h_s VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI0 mid PGATE_SL_H_N AMUXBUS_L VDDA sky130_fd_pr__pfet_g5v0d10v5 m=14 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI3 AMUXBUS_R PGATE_SR_H_N mid VDDA sky130_fd_pr__pfet_g5v0d10v5 m=14 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch_levelshifter FBK FBK_N HOLD RESET
+ SWITCH_LV SWITCH_LV_N VGND VPWR_HV VPWR_LV
*.PININFO FBK:O FBK_N:O HOLD:I RESET:I SWITCH_LV:I SWITCH_LV_N:I
*.PININFO VGND:B VPWR_HV:B VPWR_LV:B
XI184 FBK RESET VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI183 net97 VPWR_LV net109 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 FBK HOLD net105 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI182 net105 VPWR_LV net117 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net109 SWITCH_LV VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 FBK_N HOLD net97 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 net117 SWITCH_LV_N VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI185 FBK_N FBK VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 FBK FBK_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch_levelshifter

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch_s0 HOLD IN_LV OUT_H RESET VCCD VDDA
+ VSSA VSSD
*.PININFO HOLD:I IN_LV:I OUT_H:O RESET:I VCCD:B VDDA:B VSSA:B VSSD:B
XI0 net17 net13 HOLD RESET in_lv_i in_lv_n VSSA VDDA VCCD
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI22 in_lv_n IN_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 in_lv_i in_lv_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 OUT_H net13 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 in_lv_n IN_LV VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 in_lv_i in_lv_n VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 OUT_H net13 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch_s0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch_sl HOLD IN_LV OUT_H OUT_H_N RESET VCCD
+ VDDA VSSA VSSD VSWITCH
*.PININFO HOLD:I IN_LV:I OUT_H:O OUT_H_N:O RESET:I VCCD:B VDDA:B
*.PININFO VSSA:B VSSD:B VSWITCH:B
XI0 net39 net35 HOLD RESET in_lv_i in_lv_n VSSA VDDA VCCD
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI1 net48 net44 HOLD RESET in_lv_i in_lv_n VSSA VSWITCH VCCD
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI14 OUT_H net44 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 OUT_H_N net39 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 in_lv_i in_lv_n VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 in_lv_n IN_LV VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H net44 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 OUT_H_N net39 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 in_lv_i in_lv_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 in_lv_n IN_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch_sl

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amx_inv1 A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI92 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI54 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amx_inv1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat DRVHI_H DRVLO_H_N OE_H_N PD_DIS_H PU_DIS_H
+ VCC_IO VGND
*.PININFO DRVHI_H:O DRVLO_H_N:O OE_H_N:I PD_DIS_H:I PU_DIS_H:I
*.PININFO VCC_IO:I VGND:I
Xnor3_q0 oe_i_h_n DRVHI_H PD_DIS_H n1 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnor3
Xnand3_q0 oe_i_h DRVLO_H_N pu_dis_h_n n0 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe1_q0 OE_H_N oe_i_h VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_in
Xinv_oe2_q0 oe_i_h oe_i_h_n VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_in
Xinv_pudis_q0 PU_DIS_H pu_dis_h_n VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_inv_in
Xinv_out_q0 n1 DRVLO_H_N VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
Xinv_out_1_q0 n0 DRVHI_H VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
.ENDS sky130_fd_io__com_cclat

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_hvnand3 IN0 IN1 IN2 OUT VCC_IO VGND VNB
*.PININFO IN0:I IN1:I IN2:I OUT:O VCC_IO:I VGND:I VNB:I
Xmp0_q0 OUT IN0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp2_q0 OUT IN2 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp1_q0 OUT IN1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn2_q0 OUT IN2 n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn0_q0 n0 IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn1_q0 n1 IN1 n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_hvnand3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_hvnor3 IN0 IN1 IN2 OUT VCC_IO VGND VNB
*.PININFO IN0:I IN1:I IN2:I OUT:O VCC_IO:I VGND:I VNB:I
Xmp0_q0 n<0> IN0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp2_q0 OUT IN2 n<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp1_q0 n<1> IN1 n<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn0_q0 OUT IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn2_q0 OUT IN2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn1_q0 OUT IN1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_hvnor3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_i2c_fix DRVHI_H DRVLO_H_N OE_H PD_DIS_H PU_DIS_H
+ VCC_IO VGND
*.PININFO DRVHI_H:O DRVLO_H_N:O OE_H:I PD_DIS_H:I PU_DIS_H:I VCC_IO:I
*.PININFO VGND:I
Xnor3_q0 oe_i_h_n DRVHI_H PD_DIS_H n1 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnor3
Xnand3_q0 OE_H DRVLO_H_N pu_dis_h_n n0 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe2_q0 OE_H oe_i_h_n VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_in
Xinv_pudis_q0 PU_DIS_H pu_dis_h_n VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_inv_in
Xinv_out_q0 n1 DRVLO_H_N VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
Xinv_out_1_q0 n0 DRVHI_H VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
.ENDS sky130_fd_io__com_cclat_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_inv_in IN OUT VCC_IO VGND VNB
*.PININFO IN:I OUT:O VCC_IO:I VGND:I VNB:I
Xmp1_q0 OUT IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn1_q0 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_inv_in

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_inv_out IN OUT VCC_IO VGND VNB
*.PININFO IN:I OUT:O VCC_IO:I VGND:I VNB:I
XI1 OUT IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=6 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_inv_out

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_ctl_ls HLD_H_N IN OUT_H OUT_H_N RST_H SET_H VCC_IO
+ VGND VPWR
*.PININFO HLD_H_N:I IN:I OUT_H:O OUT_H_N:O RST_H:I SET_H:I VCC_IO:I
*.PININFO VGND:I VPWR:I
XI14 OUT_H_N fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 in_i in_i_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 in_i_n IN VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnset_q0 fbk_n SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 in_i in_i_n VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI58 net130 VPWR net94 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI59 net122 VPWR net98 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 fbk_n HLD_H_N net122 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI27 in_i_n IN VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 fbk HLD_H_N net130 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI3 fbk fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net98 in_i VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net94 in_i_n VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_ctl_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_inv_x1_dnw IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_inv_x1_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_nand2_dnw IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_nand2_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_nor2_dnw IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net17 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net17 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_nor2_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pad PAD VGND_IO
*.PININFO PAD:B VGND_IO:B
.ENDS sky130_fd_io__com_pad

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pddrvr_unit_2_5 ND NGIN NS
*.PININFO ND:B NGIN:I NS:B
Xndrv_q0 ND NGIN NS NS sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pddrvr_unit_2_5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pdpredrvr_pbias DRVLO_H_N EN_H EN_H_N PBIAS PD_H
+ PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_H:I EN_H_N:I PBIAS:O PD_H:I PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
XI27 n<0> PD_H EN_H_N sky130_fd_io__tk_opto
XE1 n<1> n<0> sky130_fd_io__tk_em1o
XE2 PBIAS pbias1 sky130_fd_io__tk_em1o
XE3 pbias1 net88 sky130_fd_io__tk_em1s
XE4 net108 PBIAS sky130_fd_io__tk_em1s
XE6 PBIAS net84 sky130_fd_io__tk_em1s
XE5 n<101> bias_g sky130_fd_io__tk_em1s
XI47 PBIAS bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 n<1> DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 bias_g DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 n<0> n<0> n<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 drvlo_i_h DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 bias_g n<1> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 bias_g EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 net157 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 net108 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 n<1> PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI48 n<100> PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI41 n<101> PD_H n<100> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI44 PBIAS PBIAS pbias1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 pbias1 pbias1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net183 EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net171 n<0> net183 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 PBIAS EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 drvlo_i_h DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 bias_g DRVLO_H_N net171 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 PBIAS drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 N0 VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 net161 net161 N0 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net157 net157 net161 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net88 N0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI43 net84 bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI40 N0 drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pdpredrvr_pbias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pdpredrvr_strong_slow DRVLO_H_N PD_H PDEN_H_N VCC_IO
+ VGND_IO
*.PININFO DRVLO_H_N:I PD_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
XI26 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 net25 PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 PD_H DRVLO_H_N net25 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pdpredrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pdpredrvr_weak DRVLO_H_N PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I PD_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
XI26 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 net25 PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 PD_H DRVLO_H_N net25 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pdpredrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pudrvr_strong_slow PAD PU_H_N VCC_IO VGND_IO VPB_DRVR
*.PININFO PAD:O PU_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I
Xpdrv_q0 PAD PU_H_N VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=8 w=7.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pudrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pudrvr_weak PAD PU_H_N VCC_IO VGND_IO VPB_DRVR
*.PININFO PAD:O PU_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I
Xpdrv_q0 PAD PU_H_N VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=7.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 PAD PU_H_N VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pudrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pupredrvr_nbias DRVHI_H EN_H EN_H_N NBIAS PU_H_N
+ PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_H:I EN_H_N:I NBIAS:O PU_H_N:I PUEN_H:I VCC_IO:I
*.PININFO VGND_IO:I
XI36 n<2> PU_H_N EN_H sky130_fd_io__tk_opto
XE5 NBIAS net88 sky130_fd_io__tk_em1s
XE4 n<6> net153 sky130_fd_io__tk_em1s
XE7 bias_g net90 sky130_fd_io__tk_em1s
XE6 net141 NBIAS sky130_fd_io__tk_em1s
XE1 n<2> n<1> sky130_fd_io__tk_em1o
XE2 n<6> NBIAS sky130_fd_io__tk_em1o
XI34 n<1> DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 n<1> n<2> n<2> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 bias_g n<1> VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 bias_g DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 bias_g EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 NBIAS bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 drvhi_i_h_n DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI47 n<7> bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI49 net88 bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI50 n<1> PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 VCC_IO PU_H_N net90 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 n<6> n<6> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 NBIAS NBIAS n<6> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 bias_g DRVHI_H n<3> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI27 n<3> n<2> n<4> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 n<4> EN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 drvhi_i_h_n DRVHI_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 NBIAS EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 vccio_2vtn drvhi_i_h_n VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI25 NBIAS drvhi_i_h_n VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI40 vccio_2vtn VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI39 net153 vccio_2vtn VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI44 n<8> n<8> vccio_2vtn VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI41 n<7> n<7> n<8> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI54 net141 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pupredrvr_nbias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pupredrvr_strong_slow DRVHI_H PU_H_N PUEN_H VCC_IO
+ VGND_IO
*.PININFO DRVHI_H:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XI3 PU_H_N DRVHI_H net17 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI39 net17 PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI37 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pupredrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pupredrvr_weak DRVHI_H PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XI3 PU_H_N DRVHI_H net21 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI39 net21 PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI37 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pupredrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_res_strong_slow RA RB VGND_IO
*.PININFO RA:B RB:B VGND_IO:I
XI28 net34 net30 sky130_fd_io__tk_em1s
XRI32 RB net30 sky130_fd_pr__res_generic_po W=2 L=2 m=1
XRI29 net30 net34 sky130_fd_pr__res_generic_po W=2 L=3 m=1
XRr1 net34 RA sky130_fd_pr__res_generic_po W=2 L=5 m=1
.ENDS sky130_fd_io__com_res_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_res_weak RA RB VGND_IO
*.PININFO RA:B RB:B VGND_IO:I
Xe9_q0 n<0> n<1> sky130_fd_io__tk_em1s
Xe11_q0 n<2> n<3> sky130_fd_io__tk_em1s
Xe10_q0 n<1> n<2> sky130_fd_io__tk_em1s
Xe12_q0 n<3> RB sky130_fd_io__tk_em1s
Xe13_q0 n<4> n<0> sky130_fd_io__tk_em1s
Xe14_q0 n<5> n<4> sky130_fd_io__tk_em1o
XRI84 n<0> n<1> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI62 n<3> RB sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI82 n<2> n<3> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI85 RA net64 sky130_fd_pr__res_generic_po W=0.8 L=50 m=1
XRI83 n<1> n<2> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI116 net64 n<5> sky130_fd_pr__res_generic_po W=0.8 L=12 m=1
XRI104 n<4> n<0> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
XRI134 n<5> n<4> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
.ENDS sky130_fd_io__com_res_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_xres_weak_pu RA RB VGND_IO
*.PININFO RA:B RB:B VGND_IO:I
Xe9_q0 n<0> n<1> sky130_fd_io__tk_em1s
Xe11_q0 n<2> n<3> sky130_fd_io__tk_em1s
Xe10_q0 n<1> n<2> sky130_fd_io__tk_em1s
Xe12_q0 n<3> RB sky130_fd_io__tk_em1s
Xe13_q0 n<4> n<0> sky130_fd_io__tk_em1s
Xe14_q0 n<5> n<4> sky130_fd_io__tk_em1o
XRI84 n<0> n<1> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI62 n<3> RB sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI82 n<2> n<3> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI85 RA net64 sky130_fd_pr__res_generic_po W=0.8 L=50 m=1
XRI83 n<1> n<2> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
XRI116 net64 n<5> sky130_fd_pr__res_generic_po W=0.8 L=12 m=1
XRI104 n<4> n<0> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
XRI134 n<5> n<4> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
.ENDS sky130_fd_io__com_xres_weak_pu

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__enh_nand2_1 IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__enh_nand2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__enh_nand2_1_sp IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__enh_nand2_1_sp

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__enh_nor2_x1 IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net16 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net16 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__enh_nor2_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  The local_5term cells have resistors that overlap, and the resistor
* end terminals must be added to the netlist to make it correct.

.SUBCKT sky130_fd_io__gpio_buf_localesd IN_H OUT_H OUT_VT VCC_IO VGND
+ VTRIP_SEL_H
*.PININFO IN_H:I OUT_H:O OUT_VT:O VCC_IO:B VGND:B VTRIP_SEL_H:I
Xesd_res_q0 IN_H OUT_H sky130_fd_io__res250only_small
Xggnfet2_q0 VGND OUT_VT VGND VCC_IO VGND VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet6_q0 VGND VCC_IO VGND VCC_IO OUT_H VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet5_q0 VGND VCC_IO VGND VCC_IO OUT_VT VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet1_q0 VGND OUT_H VGND VCC_IO VGND VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xhv_passgate_q0 OUT_H VTRIP_SEL_H OUT_VT VGND sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_buf_localesd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ctlv2_i2c_fix DM[2] DM[1] DM[0] DM_H[2] DM_H[1]
+ DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] ENABLE_H ENABLE_INP_H HLD_H_N HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR HYST_TRIM HYST_TRIM_H HYST_TRIM_H_N IB_MODE_SEL[1]
+ IB_MODE_SEL[0] IB_MODE_SEL_H[1] IB_MODE_SEL_H[0] IB_MODE_SEL_H_N[1]
+ IB_MODE_SEL_H_N[0] INP_DIS INP_DIS_H_N OD_I_H_N SLEW_CTL[1] SLEW_CTL[0]
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] VCCD VDDIO_Q VSSD
+ VTRIP_SEL VTRIP_SEL_H
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O ENABLE_H:I
*.PININFO ENABLE_INP_H:I HLD_H_N:I HLD_I_H_N:O HLD_I_OVR_H:O HLD_OVR:I
*.PININFO HYST_TRIM:I HYST_TRIM_H:O HYST_TRIM_H_N:O IB_MODE_SEL[1]:I
*.PININFO IB_MODE_SEL[0]:I IB_MODE_SEL_H[1]:O IB_MODE_SEL_H[0]:O
*.PININFO IB_MODE_SEL_H_N[1]:O IB_MODE_SEL_H_N[0]:O INP_DIS:I
*.PININFO INP_DIS_H_N:O OD_I_H_N:O SLEW_CTL[1]:I SLEW_CTL[0]:I
*.PININFO SLEW_CTL_H[1]:O SLEW_CTL_H[0]:O SLEW_CTL_H_N[1]:O
*.PININFO SLEW_CTL_H_N[0]:O VCCD:I VDDIO_Q:I VSSD:I VTRIP_SEL:I
*.PININFO VTRIP_SEL_H:O
Xls_bank_q0 DM[2] DM[1] DM[0] DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N HYST_TRIM HYST_TRIM_H HYST_TRIM_H_N IB_MODE_SEL[1]
+ IB_MODE_SEL[0] IB_MODE_SEL_H[1] IB_MODE_SEL_H[0] IB_MODE_SEL_H_N[1]
+ IB_MODE_SEL_H_N[0] INP_DIS net83 INP_DIS_H_N OD_I_H_N SLEW_CTL[1] SLEW_CTL[0]
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] startup_rst_h
+ inp_startup_en_h VDDIO_Q VSSD VCCD VTRIP_SEL VTRIP_SEL_H net77
+ sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix
Xhld_dis_blk_q0 ENABLE_H HLD_H_N HLD_I_H_N HLD_I_OVR_H HLD_OVR OD_I_H_N VDDIO_Q
+ VSSD VCCD sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix
XI75 ENABLE_INP_H ENABLE_H startup_rst_h VSSD VDDIO_Q sky130_fd_io__hvsbt_nor
XI56 net109 ENABLE_INP_H net108 VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI77 OD_I_H_N net109 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI57 net108 inp_startup_en_h VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpio_ctlv2_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_dat_ls HLD_H_N IN OUT_H OUT_H_N RST_H SET_H VCC_IO
+ VGND VPWR_KA
*.PININFO HLD_H_N:I IN:I OUT_H:O OUT_H_N:O RST_H:I SET_H:I VCC_IO:I
*.PININFO VGND:I VPWR_KA:I
XI3 fbk fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 fbk HLD_H_N net79 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 fbk_n HLD_H_N net83 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net107 in_i_n VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net103 in_i VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnset_q0 fbk_n SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 in_i_n IN VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 in_i in_i_n VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net83 VPWR_KA net103 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net79 VPWR_KA net107 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 in_i in_i_n VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 OUT_H_N fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 in_i_n IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_dat_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_dat_ls_i2c_fix HLD_H_N IN OUT_H_N SET_H SET_H_N
+ VCC_IO VGND VPWR_KA
*.PININFO HLD_H_N:I IN:I OUT_H_N:O SET_H:I SET_H_N:I VCC_IO:I VGND:I
*.PININFO VPWR_KA:I
XI3 fbk fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 fbk HLD_H_N net76 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 fbk_n HLD_H_N net80 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net100 in_i_n VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net96 in_i VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnset_q0 fbk_n SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 in_i_n IN VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 in_i in_i_n VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net80 VPWR_KA net96 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net76 VPWR_KA net100 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 in_i in_i_n VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 OUT_H_N fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 fbk SET_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 in_i_n IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_dat_ls_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_amux_i2c_fix AMUXBUS_A AMUXBUS_B ANALOG_EN
+ ANALOG_POL ANALOG_SEL ENABLE_VDDA_H ENABLE_VSWITCH_H HLD_I_H_N NGA_PAD_VPMP_H
+ NGB_PAD_VPMP_H NGHS_H OUT PAD PD_CSD_H PGHS_H PU_CSD_H PUG_H[1] PUG_H[0] VCCD
+ VDDA VDDIO VDDIO_Q VPB_DRVR VSSA VSSD VSSIO VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I ENABLE_VDDA_H:I ENABLE_VSWITCH_H:I HLD_I_H_N:I
*.PININFO NGA_PAD_VPMP_H:O NGB_PAD_VPMP_H:O NGHS_H:I OUT:I PAD:B
*.PININFO PD_CSD_H:O PGHS_H:I PU_CSD_H:O PUG_H[1]:B PUG_H[0]:B VCCD:I
*.PININFO VDDA:I VDDIO:I VDDIO_Q:I VPB_DRVR:B VSSA:I VSSD:I VSSIO:I
*.PININFO VSWITCH:I
XI78 HLD_I_H_N hld_i_h_amux_sw VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XBBM_logic ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H enable_vdda_h_n
+ ENABLE_VSWITCH_H HLD_I_H_N nga_amx_vpmp_h NGA_PAD_VPMP_H ngb_amx_vpmp_h
+ NGB_PAD_VPMP_H nmida_vccd nmidb_vccd OUT PD_CSD_H pga_amx_vdda_h_n
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n PU_CSD_H VCCD VDDA
+ VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix
xI77 VSSA VDDA sky130_fd_io__condiode
XI26 net128 net142 sky130_fd_io__res75only_small
XI58 net126 net139 sky130_fd_io__res75only_small
XI28 net124 net144 sky130_fd_io__res75only_small
XI57 PAD net126 sky130_fd_io__res75only_small
XI27 net120 net143 sky130_fd_io__res75only_small
XI55 PAD net128 sky130_fd_io__res75only_small
XI54 PAD net124 sky130_fd_io__res75only_small
XI53 PAD net120 sky130_fd_io__res75only_small
Xmux_a_q0 AMUXBUS_A nga_amx_vpmp_h NGA_PAD_VPMP_H NGHS_H nmida_vccd net144
+ net144 net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n PGHS_H PUG_H[0] VDDA VDDIO VPB_DRVR VSSA
+ VSSD VSSIO sky130_fd_io__gpio_ovtv2_amux_switch
Xmux_b_q0 AMUXBUS_B ngb_amx_vpmp_h NGB_PAD_VPMP_H NGHS_H nmidb_vccd net144
+ net144 net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw
+ pgb_amx_vdda_h_n pgb_pad_vddioq_h_n PGHS_H PUG_H[1] VDDA VDDIO VPB_DRVR VSSA
+ VSSD VSSIO sky130_fd_io__gpio_ovtv2_amux_switch
.ENDS sky130_fd_io__gpio_ovtv2_amux_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_amux_switch AG_HV NG_AG_VPMP NG_PAD_VPMP NGHS_H
+ NMID_VDDA PAD_HV_N0 PAD_HV_N1 PAD_HV_N2 PAD_HV_N3 PAD_HV_P0 PAD_HV_P1 PD_H_VDDA
+ PD_H_VDDIO PG_AG_VDDA PG_PAD_VDDIOQ PGHS_H PUG_H VDDA VDDIO VPB_DRVR VSSA VSSD
+ VSSIO
*.PININFO AG_HV:B NG_AG_VPMP:I NG_PAD_VPMP:I NGHS_H:I NMID_VDDA:I
*.PININFO PAD_HV_N0:B PAD_HV_N1:B PAD_HV_N2:B PAD_HV_N3:B PAD_HV_P0:B
*.PININFO PAD_HV_P1:B PD_H_VDDA:I PD_H_VDDIO:I PG_AG_VDDA:I
*.PININFO PG_PAD_VDDIOQ:I PGHS_H:I PUG_H:B VDDA:I VDDIO:I VPB_DRVR:B
*.PININFO VSSA:I VSSD:I VSSIO:I
xI72 VSSA VDDIO sky130_fd_io__condiode
xI71 mid1 VDDIO sky130_fd_io__condiode
xI70 mid VDDIO sky130_fd_io__condiode
XI56 VSSA net85 sky130_fd_io__res75only_small
XI12 VSSA net83 sky130_fd_io__res75only_small
XI46 PAD_HV_N3 NG_PAD_VPMP mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 mid NG_PAD_VPMP PAD_HV_N1 mid sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 PAD_HV_N0 NG_PAD_VPMP mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 mid1 NG_PAD_VPMP PAD_HV_N2 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 mid NG_AG_VPMP AG_HV mid sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI57 mid1 NMID_VDDA net85 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI63 PUG_H NGHS_H PG_PAD_VDDIOQ VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI47 mid1 NG_AG_VPMP AG_HV mid1 sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI75<1> mid PD_H_VDDA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI75<0> mid1 PD_H_VDDA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74<1> mid PD_H_VDDIO VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74<0> mid1 PD_H_VDDIO VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 mid NMID_VDDA net83 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 mid PUG_H PAD_HV_P1 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 mid PUG_H PAD_HV_P0 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI62 PG_PAD_VDDIOQ PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 mid PG_AG_VDDA AG_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 m=4 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_amux_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim to add the additional pin on signal_5_sym_hv_local_5term
* needed to represent the connection from the end of the annular m1 resistor
* (short) back to VDDIO_Q

.SUBCKT sky130_fd_io__gpio_ovtv2_buf_localesd IN_H OUT_H OUT_VT VDDIO_Q VSSD
+ VTRIP_SEL_H
*.PININFO IN_H:I OUT_H:O OUT_VT:O VDDIO_Q:B VSSD:B VTRIP_SEL_H:I
Xesd_res_q0 IN_H OUT_H sky130_fd_io__res250only_small
Xggnfet6_q0 VSSD VDDIO_Q VSSD VDDIO_Q OUT_H noconnect1
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet1_q0 VSSD OUT_H VSSD VDDIO_Q VSSD noconnect2
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xhv_passgate_q0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_buf_localesd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix ENABLE_H HLD_H_N HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR OD_I_H_N VCC_IO VGND VPWR
*.PININFO ENABLE_H:I HLD_H_N:I HLD_I_H_N:O HLD_I_OVR_H:O HLD_OVR:I
*.PININFO OD_I_H_N:O VCC_IO:I VGND:I VPWR:I
Xhld_nand_q0 ENABLE_H HLD_H_N n1 VGND VCC_IO sky130_fd_io__enh_nand2_1_sp
XI50 OD_I_H_N net45 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI46 n1 n1 n2 VGND VCC_IO sky130_fd_io__enh_nor2_x1
XI49 od_h od_h OD_I_H_N VGND VCC_IO sky130_fd_io__enh_nor2_x1
XI48 ENABLE_H ENABLE_H od_h VGND VCC_IO sky130_fd_io__enh_nand2_1
XI155 n3 n3 HLD_I_H_N VGND VCC_IO sky130_fd_io__nor2_4_enhpath
XI154 n2 n2 n3 VGND VCC_IO sky130_fd_io__nand2_2_enhpath
Xhld_ovr_ls_q0 n2 HLD_OVR hld_ovr_h net79 od_h VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
XI30 net45 hld_i_ovr_h_n HLD_I_OVR_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI26 n2 hld_ovr_h hld_i_ovr_h_n VGND VCC_IO sky130_fd_io__hvsbt_nor
.ENDS sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix DM[2] DM[1] DM[0] DM_H[2]
+ DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N HYST_TRIM HYST_TRIM_H
+ HYST_TRIM_H_N IB_MODE_SEL[1] IB_MODE_SEL[0] IB_MODE_SEL_H[1] IB_MODE_SEL_H[0]
+ IB_MODE_SEL_H_N[1] IB_MODE_SEL_H_N[0] INP_DIS INP_DIS_H INP_DIS_H_N OD_I_H_N
+ SLEW_CTL[1] SLEW_CTL[0] SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1]
+ SLEW_CTL_H_N[0] STARTUP_RST_H STARTUP_ST_H VCC_IO VGND VPWR VTRIP_SEL
+ VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O HLD_I_H_N:I HYST_TRIM:I
*.PININFO HYST_TRIM_H:O HYST_TRIM_H_N:O IB_MODE_SEL[1]:I
*.PININFO IB_MODE_SEL[0]:I IB_MODE_SEL_H[1]:O IB_MODE_SEL_H[0]:O
*.PININFO IB_MODE_SEL_H_N[1]:O IB_MODE_SEL_H_N[0]:O INP_DIS:I
*.PININFO INP_DIS_H:O INP_DIS_H_N:O OD_I_H_N:I SLEW_CTL[1]:I
*.PININFO SLEW_CTL[0]:I SLEW_CTL_H[1]:O SLEW_CTL_H[0]:O
*.PININFO SLEW_CTL_H_N[1]:O SLEW_CTL_H_N[0]:O STARTUP_RST_H:I
*.PININFO STARTUP_ST_H:I VCC_IO:I VGND:I VPWR:I VTRIP_SEL:I
*.PININFO VTRIP_SEL_H:O VTRIP_SEL_H_N:O
XI836 OD_I_H_N od_i_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
Xtrip_sel_st_q0 trip_sel_st_h od_i_h VGND sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> od_i_h VGND sky130_fd_io__tk_optiA
Xtrip_sel_rst_q0 trip_sel_rst_h VGND od_i_h sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> od_i_h VGND sky130_fd_io__tk_optiA
XI804<1> dm_rst_h<2> VGND od_i_h sky130_fd_io__tk_optiC
XI338<1> dm_rst_h<0> STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_optiC
XI615 hyst_trim_st_h od_i_h VGND sky130_fd_io__tk_opti
XI614 hyst_trim_rst_h VGND od_i_h sky130_fd_io__tk_opti
XI598<1> ib_mode_sel_st_h<1> od_i_h VGND sky130_fd_io__tk_opti
XI598<0> ib_mode_sel_st_h<0> od_i_h VGND sky130_fd_io__tk_opti
XI597<1> ib_mode_sel_rst_h<1> VGND od_i_h sky130_fd_io__tk_opti
XI597<0> ib_mode_sel_rst_h<0> VGND od_i_h sky130_fd_io__tk_opti
XI337<1> dm_st_h<0> STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_optiA
XI805<1> dm_rst_h<1> VGND od_i_h sky130_fd_io__tk_optiC
XI666<1> slew_ctl_st_h<1> od_i_h VGND sky130_fd_io__tk_opti
XI666<0> slew_ctl_st_h<0> od_i_h VGND sky130_fd_io__tk_opti
XI665<1> slew_ctl_rst_h<1> VGND od_i_h sky130_fd_io__tk_opti
XI665<0> slew_ctl_rst_h<0> VGND od_i_h sky130_fd_io__tk_opti
XI687 ie_n_st_h STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_optiC
XI686 ie_n_rst_h STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_optiA
Xdm_ls_0_q0 HLD_I_H_N DM[0] DM_H[0] DM_H_N[0] dm_rst_h<0> dm_st_h<0> VCC_IO VGND
+ VPWR sky130_fd_io__com_ctl_ls
Xinp_dis_ls_q0 HLD_I_H_N INP_DIS INP_DIS_H INP_DIS_H_N ie_n_rst_h ie_n_st_h
+ VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xtrip_sel_ls_q0 HLD_I_H_N VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N trip_sel_rst_h
+ trip_sel_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
XI616 HLD_I_H_N HYST_TRIM HYST_TRIM_H HYST_TRIM_H_N hyst_trim_rst_h
+ hyst_trim_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
XI595<1> HLD_I_H_N IB_MODE_SEL[1] IB_MODE_SEL_H[1] IB_MODE_SEL_H_N[1]
+ ib_mode_sel_rst_h<1> ib_mode_sel_st_h<1> VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
XI595<0> HLD_I_H_N IB_MODE_SEL[0] IB_MODE_SEL_H[0] IB_MODE_SEL_H_N[0]
+ ib_mode_sel_rst_h<0> ib_mode_sel_st_h<0> VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
XI667<1> HLD_I_H_N SLEW_CTL[1] SLEW_CTL_H[1] SLEW_CTL_H_N[1] slew_ctl_rst_h<1>
+ slew_ctl_st_h<1> VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
XI667<0> HLD_I_H_N SLEW_CTL[0] SLEW_CTL_H[0] SLEW_CTL_H_N[0] slew_ctl_rst_h<0>
+ slew_ctl_st_h<0> VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<2>_q0 HLD_I_H_N DM[2] DM_H[2] DM_H_N[2] dm_rst_h<2> dm_st_h<2> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<1>_q0 HLD_I_H_N DM[1] DM_H[1] DM_H_N[1] dm_rst_h<1> dm_st_h<1> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_bias PSWG_H VCC_IO VPB_DRVR
*.PININFO PSWG_H:I VCC_IO:I VPB_DRVR:O
Xpsw_vccio_q0 VPB_DRVR PSWG_H VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=22
+ w=15.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI36 VPB_DRVR PSWG_H VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=9 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_bias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix EN_H ENHS_LAT_H_N
+ FORCEHI_H[1] OD_I_H_N P3OUT PAD_ESD PGHS_H VDDIO VPB_DRVR VPWR_KA VSSD
*.PININFO EN_H:I ENHS_LAT_H_N:O FORCEHI_H[1]:I OD_I_H_N:I P3OUT:O
*.PININFO PAD_ESD:I PGHS_H:B VDDIO:I VPB_DRVR:I VPWR_KA:I VSSD:I
Xhslog_q0 dishs_h dishs_h_n EN_H enhs_h enhs_h_n enhs_lathys_h_n exiths_h
+ FORCEHI_H[1] OD_I_H_N VDDIO VSSD sky130_fd_io__sio_hotswap_log_i2c_fix
Xhslatch_q0 dishs_h dishs_h_n enhs_h enhs_h_n ENHS_LAT_H_N enhs_lathys_h_n
+ exiths_h P3OUT PAD_ESD PGHS_H VDDIO VSSD VPB_DRVR VPWR_KA
+ sky130_fd_io__gpio_ovtv2_hotswap_latch
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix FORCE_H[1] NGHS_H
+ OD_I_H_N OE_HS_H P2G PAD PAD_ESD PGHS_H PUG_H[7] PUG_H[6] PUG_H[5] PUG_H[4]
+ PUG_H[3] PUG_H[2] PUG_H[1] PUG_H[0] VCC_IO_SOFT VDDIO VPB_DRVR VPWR_KA VSSD
*.PININFO FORCE_H[1]:I NGHS_H:O OD_I_H_N:I OE_HS_H:I P2G:O PAD:I
*.PININFO PAD_ESD:I PGHS_H:O PUG_H[7]:B PUG_H[6]:B PUG_H[5]:B
*.PININFO PUG_H[4]:B PUG_H[3]:B PUG_H[2]:B PUG_H[1]:B PUG_H[0]:B
*.PININFO VCC_IO_SOFT:O VDDIO:I VPB_DRVR:O VPWR_KA:I VSSD:I
Xnon_overlap_q0 p1g NGHS_H P2G padlo VSSD VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix
Xpug47_q0 padlo PUG_H[4] PUG_H[7] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix
Xpghs_q0 OE_HS_H FORCE_H[1] OD_I_H_N net74 PAD_ESD padlo p1g tie_hi VCC_IO_SOFT
+ VDDIO VPB_DRVR VPWR_KA VSSD sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix
Xresd_tiehi_q0 VPB_DRVR tie_hi sky130_fd_io__sio_tk_tie_r_out_esd
Xresd_vccio_q0 VDDIO VCC_IO_SOFT sky130_fd_io__sio_tk_tie_r_out_esd
Xpug<3>_q0 PAD_ESD padlo PUG_H[3] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<2>_q0 PAD_ESD padlo PUG_H[2] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<1>_q0 PAD_ESD padlo PUG_H[1] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<0>_q0 PAD_ESD padlo PUG_H[0] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<6>_q0 PAD_ESD padlo PUG_H[6] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<5>_q0 PAD_ESD padlo PUG_H[5] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xp1_bias_q0 p1g VDDIO VPB_DRVR sky130_fd_io__gpio_ovtv2_hotswap_bias
Xp2p4_bias_q0 P2G PAD VCC_IO_SOFT VCC_IO_SOFT VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias
* RI26 P2G net137 short
* RI39 P2G net74 short
* RI49 PGHS_H p1g short
RI26 P2G net137 sky130_fd_pr__res_generic_m1 W=0.4 L=0.01
RI39 P2G net74 sky130_fd_pr__res_generic_m1 W=0.4 L=0.01
RI49 PGHS_H p1g sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_latch DISHS_H DISHS_H_N ENHS_H ENHS_H_N
+ ENHS_LAT_H_N ENHS_LATHYS_H_N EXITHS_H P3OUT PAD_ESD PGHS_H VCC_IO VGND VPB_DRVR
+ VPWR_KA
*.PININFO DISHS_H:I DISHS_H_N:I ENHS_H:I ENHS_H_N:I ENHS_LAT_H_N:O
*.PININFO ENHS_LATHYS_H_N:O EXITHS_H:I P3OUT:O PAD_ESD:I PGHS_H:B
*.PININFO VCC_IO:I VGND:I VPB_DRVR:I VPWR_KA:I
XI660 VGND net102 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI528 n6 net96 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XEhys2 ENHS_LATHYS_H_N ENHS_LAT_H_N sky130_fd_io__tk_em1o
XI658 net96 ENHS_LAT_H_N sky130_fd_io__tk_em1s
XEhys1 net117 ENHS_LATHYS_H_N sky130_fd_io__tk_em1s
Xhys_q0 n6 net117 VCC_IO VGND sky130_fd_io__sio_hotswap_hys
Xpghspd_q0 ENHS_H n2 PGHS_H VGND sky130_fd_io__sio_hotswap_pghspd
Xwpdenhs_q0 VPWR_KA net127 VGND sky130_fd_io__sio_hotswap_wpd
Xwpdexhs_q0 VPWR_KA net124 VGND sky130_fd_io__sio_hotswap_wpd
XI502 net186 PGHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI484 net161 ENHS_H PGHS_H VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI491 n5 n6 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI498 n2 n6 net124 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI500 net170 ENHS_H_N n2 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnexiths_q0 PGHS_H EXITHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI485 n3 n2 net161 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI499 n4 PGHS_H net170 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI497 n6 n5 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xndishs_q0 PGHS_H DISHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI508 n2 ENHS_H_N net186 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI696 VGND EXITHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI487 PGHS_H n5 net127 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI697 VGND DISHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI492 n5 n6 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI503 n4 VGND VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI488 n3 VGND VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI505 n6 n5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI493 n5 n3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI323 n2 DISHS_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI279 n2 PAD_ESD VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI504 n6 n4 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI689 P3OUT PAD_ESD VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=12 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_latch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix P1G P1GB P2G PADLO
+ VGND VPWR
*.PININFO P1G:O P1GB:O P2G:O PADLO:I VGND:I VPWR:I
XI76 P1G P1GB VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI64 p1g_new PADLO VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 padlo_bar PADLO VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI50 p2g_new p1g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI49 p2g_new padlo_bar VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI65 p1g_new p2g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77 P2G p2gb VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI70 p2gb p2g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI72 P1GB p1g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI54 padlo_bar PADLO VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI69 p1g_new PADLO net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI78 P2G p2gb VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI67 net140 p2g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI71 p2gb p2g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI79 P1G P1GB VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI51 p2g_new padlo_bar net124 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI73 P1GB p1g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI52 net124 p1g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix EN_H FORCE_H[1] OD_I_H_N
+ P3OUT PAD PADLO PGHS_H TIE_HI VCC_IO_SOFT VDDIO VPB_DRVR VPWR_KA VSSD
*.PININFO EN_H:I FORCE_H[1]:I OD_I_H_N:I P3OUT:O PAD:I PADLO:O
*.PININFO PGHS_H:O TIE_HI:I VCC_IO_SOFT:I VDDIO:I VPB_DRVR:I VPWR_KA:I
*.PININFO VSSD:I
Xhsctl_q0 EN_H enhs_lat_h_n FORCE_H[1] OD_I_H_N P3OUT PAD net50 VDDIO VPB_DRVR
+ VPWR_KA VSSD sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix
XI3 enhs_latbuf_h_n PADLO sky130_fd_io__sio_tk_em1s
XEpghs12 PGHS_H net54 sky130_fd_io__sio_tk_em1o
XI2 enhs_lat_h enhs_latbuf_h_n VSSD VSSD VDDIO VDDIO
+ sky130_fd_io__gpio_ovtv2_hvsbt_inv_x4
XI1 enhs_lat_h_n enhs_lat_h VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x1
Xpghspu_q0 PAD PGHS_H net50 TIE_HI VCC_IO_SOFT VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pghspu
Xclamp_q0 VSSD VDDIO VSSD VDDIO PAD noconnect sky130_fd_io__signal_5_sym_hv_local_5term
Xpghs12_q0 net54 PADLO VPB_DRVR VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0
+ l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghspu PAD PGHS_H PGHS_H_LATCH TIE_HI
+ VCC_IO_SOFT VPB_DRVR
*.PININFO PAD:I PGHS_H:O PGHS_H_LATCH:O TIE_HI:I VCC_IO_SOFT:I
*.PININFO VPB_DRVR:I
XEg9 TIE_HI pg8 sky130_fd_io__sio_tk_em1o
XEg2 pg2 VCC_IO_SOFT sky130_fd_io__sio_tk_em1s
XEg5 pg6 pg4 sky130_fd_io__sio_tk_em1s
XEg4 pg4 pg3 sky130_fd_io__sio_tk_em1s
XEpghs3 padhi3 PGHS_H_LATCH sky130_fd_io__sio_tk_em1s
XEg3 pg3 pg2 sky130_fd_io__sio_tk_em1s
XEpghs7 padhi7 net36 sky130_fd_io__sio_tk_em1s
XEg7 pg7 pg6 sky130_fd_io__sio_tk_em1s
XEg8 pg8 pg7 sky130_fd_io__sio_tk_em1s
XEpghs2 padhi2 padhi3 sky130_fd_io__sio_tk_em1s
XEpghs8 PGHS_H padhi7 sky130_fd_io__sio_tk_em1s
Xpghs8_q0 PGHS_H pg8 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs2_q0 padhi2 pg2 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs3_q0 padhi3 pg3 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs6_q0 net36 pg6 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs4_q0 PGHS_H_LATCH pg4 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs7_q0 padhi7 pg7 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pghspu

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug PAD PADLO PUG_H TIE_HI VPB_DRVR
*.PININFO PAD:I PADLO:I PUG_H:O TIE_HI:I VPB_DRVR:I
XEg1 PADLO net22 sky130_fd_io__sio_tk_em1s
XI65 net24 TIE_HI sky130_fd_io__sio_tk_em2s
XEs2 net26 TIE_HI sky130_fd_io__sio_tk_em2s
XEs1 PAD net26 sky130_fd_io__sio_tk_em2o
XEg2 net22 net24 sky130_fd_io__sio_tk_em2o
XI52 PUG_H net22 net26 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=1.825 sb=1.825 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 PUG_H net24 net26 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pug

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix PADLO PUG4_H PUG7_H TIE_HI
+ VPB_DRVR
*.PININFO PADLO:I PUG4_H:O PUG7_H:O TIE_HI:I VPB_DRVR:I
XI52 PUG4_H PADLO TIE_HI VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=1.825 sb=1.825 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 PUG7_H PADLO TIE_HI VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias P2G PAD SOFT_VCC_IO TIE_HI
+ VPB_DRVR
*.PININFO P2G:I PAD:I SOFT_VCC_IO:I TIE_HI:I VPB_DRVR:B
Xpsw_pad4_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad0_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad3_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad2_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad5_q0 VPB_DRVR VPB_DRVR SOFT_VCC_IO PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad1_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
XI5 TIE_HI SOFT_VCC_IO sky130_fd_io__tk_em2o
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit PB PD PGIN PS
*.PININFO PB:I PD:B PGIN:I PS:B
Xpdrv_q0 PD PGIN PS PB sky130_fd_pr__esd_pfet_g5v0d10v5 m=2 w=15.5 l=0.55 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ibuf_se EN_H EN_H_N ENABLE_VDDIO_LV IBUFMUX_OUT
+ IBUFMUX_OUT_H IN_H IN_VT MODE_NORMAL_N MODE_REF_3V_N MODE_REF_N MODE_VCCD_N
+ VCCHIB VDDIO_Q VREFIN VSSD VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO EN_H:I EN_H_N:I ENABLE_VDDIO_LV:I IBUFMUX_OUT:O
*.PININFO IBUFMUX_OUT_H:O IN_H:I IN_VT:I MODE_NORMAL_N:I
*.PININFO MODE_REF_3V_N:I MODE_REF_N:I MODE_VCCD_N:I VCCHIB:I
*.PININFO VDDIO_Q:I VREFIN:I VSSD:I VTRIP_SEL_H:I VTRIP_SEL_H_N:I
Xlvls_q0 ENABLE_VDDIO_LV out IBUFMUX_OUT net43 VCCHIB VSSD
+ sky130_fd_io__gpio_ovtv2_ipath_lvls
Xhvls_q0 EN_H_N out out_n IBUFMUX_OUT_H net49 VDDIO_Q VSSD
+ sky130_fd_io__gpio_ovtv2_ipath_hvls
Xbuf_q0 EN_H EN_H_N ENABLE_VDDIO_LV IN_H IN_VT MODE_NORMAL_N MODE_REF_3V_N
+ MODE_REF_N MODE_VCCD_N out out_n VCCHIB VDDIO_Q VREFIN VSSD VTRIP_SEL_H
+ VTRIP_SEL_H_N sky130_fd_io__gpio_ovtv2_in_buf
.ENDS sky130_fd_io__gpio_ovtv2_ibuf_se

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ictl_logic DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ HYS_TRIM IBUF_MODE_SEL[0] IBUF_MODE_SEL[1] INP_DIS_H_N INP_DIS_I_H INP_DIS_I_H_N
+ MODE_NORMAL_N MODE_REF_3V_N MODE_REF_N MODE_VCCD_N TRIPSEL_I_H TRIPSEL_I_H_N
+ VDDIO_Q VSSD VTRIP_SEL_H
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I HYS_TRIM:I
*.PININFO IBUF_MODE_SEL[0]:I IBUF_MODE_SEL[1]:I INP_DIS_H_N:I
*.PININFO INP_DIS_I_H:O INP_DIS_I_H_N:O MODE_NORMAL_N:O
*.PININFO MODE_REF_3V_N:O MODE_REF_N:O MODE_VCCD_N:O TRIPSEL_I_H:O
*.PININFO TRIPSEL_I_H_N:O VDDIO_Q:I VSSD:I VTRIP_SEL_H:I
XI41 net66 MODE_NORMAL_N TRIPSEL_I_H VSSD VDDIO_Q sky130_fd_io__hvsbt_nor
XI34 IBUF_MODE_SEL[1] net70 net60 VSSD VDDIO_Q sky130_fd_io__hvsbt_nor
XI33 IBUF_MODE_SEL[1] IBUF_MODE_SEL[0] net55 VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
Xdm10nand_inv_q0 nand_dm01 and_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI68 INP_DIS_I_H INP_DIS_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI43 TRIPSEL_I_H TRIPSEL_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI50 MODE_REF_N mode_ref VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI39 IBUF_MODE_SEL[0] net70 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI61 VTRIP_SEL_H net66 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
Xinpdis_q0 dm_buf_dis INP_DIS_H_N INP_DIS_I_H VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
Xdm210_q0 DM_H_N[2] and_dm01 dm_buf_dis VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
Xdm10_q0 DM_H_N[1] DM_H_N[0] nand_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI40 INP_DIS_I_H_N IBUF_MODE_SEL[1] MODE_REF_N VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
XI36 INP_DIS_I_H_N net60 MODE_VCCD_N VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI35 INP_DIS_I_H_N net55 MODE_NORMAL_N VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI52 mode_ref HYS_TRIM MODE_REF_3V_N VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
.ENDS sky130_fd_io__gpio_ovtv2_ictl_logic

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_in_buf EN_H EN_H_N ENABLE_VDDIO_LV IN_H IN_VT
+ MODE_NORMAL_N MODE_REF_3V_N MODE_REF_N MODE_VCCD_N OUT OUT_N VCCHIB VDDIO_Q
+ VREFIN VSSD VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO EN_H:I EN_H_N:I ENABLE_VDDIO_LV:I IN_H:I IN_VT:I
*.PININFO MODE_NORMAL_N:I MODE_REF_3V_N:I MODE_REF_N:I MODE_VCCD_N:I
*.PININFO OUT:O OUT_N:O VCCHIB:I VDDIO_Q:I VREFIN:I VSSD:I
*.PININFO VTRIP_SEL_H:I VTRIP_SEL_H_N:I
XI35 ENABLE_VDDIO_LV EN_H enable_vddio_lv_n VSSD VCCHIB
+ sky130_fd_io__hvsbt_nand2
xI405 virt_pwr1 VDDIO_Q sky130_fd_io__condiode
xI404 virt_pwr VDDIO_Q sky130_fd_io__condiode
XI488 VTRIP_SEL_H MODE_NORMAL_N mode_normal_cmos_h VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
XI43 mode_normal_cmos_h mode_normal_cmos_h_n VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_inv_x1
XI630 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI105 fbk1 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI620 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI441 IN_VT VTRIP_SEL_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI417 OUT EN_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI419 OUT_N EN_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI394 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI494 fbk IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 fbk2 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 OUT in_b VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI49 vddio_ref VREFIN virt_pwr virt_pwr sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0
+ l=0.9 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI451 fbk IN_VT VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=12 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI453 in_b IN_H fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI111 vddio_ref1 VREFIN virt_pwr1 virt_pwr1 sky130_fd_pr__nfet_05v0_nvt m=3
+ w=10.0 l=0.9 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI446 OUT_N OUT VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI389 virt_pwr VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI450 in_b IN_VT fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI274 fbk1 MODE_REF_N virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI116 virt_pwr MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI109 in_b IN_H virt_pwr virt_pwr sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT in_b virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 fbk2 mode_normal_cmos_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI611 fbk1 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI396 vddio_ref1 MODE_REF_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI115 virt_pwr MODE_VCCD_N vcchib_int virt_pwr sky130_fd_pr__pfet_g5v0d10v5 m=4
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI478 vcchib_int1 enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=8
+ w=5.0 l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI373 vddio_ref MODE_REF_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI403 OUT in_b virt_pwr2 virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI376 fbk2 MODE_REF_3V_N virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=4
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI477 vcchib_int enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=8
+ w=5.0 l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI401 in_b IN_H virt_pwr2 virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI457 OUT_N OUT virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI486 fbk1 MODE_VCCD_N vcchib_int virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI400 virt_pwr2 MODE_VCCD_N vcchib_int virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI381 virt_pwr1 MODE_VCCD_N vcchib_int1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5
+ m=6 w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI380 virt_pwr1 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ipath DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ ENABLE_VDDIO_LV HYS_TRIM_H IB_MODE_SEL_H[1] IB_MODE_SEL_H[0] INP_DIS_H_N OUT
+ OUT_H PAD VCCHIB VDDIO_Q VINREF VSSD VTRIP_SEL_H
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I ENABLE_VDDIO_LV:I
*.PININFO HYS_TRIM_H:I IB_MODE_SEL_H[1]:I IB_MODE_SEL_H[0]:I
*.PININFO INP_DIS_H_N:I OUT:O OUT_H:O PAD:B VCCHIB:I VDDIO_Q:I
*.PININFO VINREF:B VSSD:I VTRIP_SEL_H:I
Xibuf_se_q0 en_h en_h_n ENABLE_VDDIO_LV OUT OUT_H in_h in_vt mode_normal_n
+ mode_ref_3v_n mode_ref_n mode_vccd_n VCCHIB VDDIO_Q VINREF VSSD tripsel_i_h
+ tripsel_i_h_n sky130_fd_io__gpio_ovtv2_ibuf_se
Xesd_q0 PAD in_h in_vt VDDIO_Q VSSD tripsel_i_h
+ sky130_fd_io__gpio_ovtv2_buf_localesd
Xlogic_q0 DM_H_N[2] DM_H_N[1] DM_H_N[0] HYS_TRIM_H IB_MODE_SEL_H[0]
+ IB_MODE_SEL_H[1] INP_DIS_H_N en_h_n en_h mode_normal_n mode_ref_3v_n mode_ref_n
+ mode_vccd_n tripsel_i_h tripsel_i_h_n VDDIO_Q VSSD VTRIP_SEL_H
+ sky130_fd_io__gpio_ovtv2_ictl_logic
.ENDS sky130_fd_io__gpio_ovtv2_ipath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_hvls EN_H_N IN INB OUT OUT_B VDDIO_Q VSSD
*.PININFO EN_H_N:I IN:I INB:I OUT:O OUT_B:O VDDIO_Q:I VSSD:I
XI250 fbk fbk_b VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI253 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI249 fbk_b fbk VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248 OUT_B fbk VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI247 OUT_B fbk VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI252 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI304 fbk INB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI262 fbk EN_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI246 fbk_b IN VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_ipath_hvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_lvls ENABLE_VDDIO_LV IN OUT OUT_B VCCHIB
+ VSSD
*.PININFO ENABLE_VDDIO_LV:I IN:I OUT:O OUT_B:O VCCHIB:I VSSD:I
XI248 fbk_n IN VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI271 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8_hvt m=2 w=5.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI281 fbk_n ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI272 OUT_B fbk VCCHIB VCCHIB sky130_fd_pr__pfet_01v8_hvt m=1 w=5.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI277 fbk fbk_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8_hvt m=1 w=5.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI273 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI278 fbk fbk_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI305 OUT_B fbk VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI535 fbk_n IN vssd_1 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI279 vssd_1 ENABLE_VDDIO_LV VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_ipath_lvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix DRVHI_H DRVLO_H_N
+ I2C_MODE_H_N NGHS_H OE_I_H_N PAD PD_DIS_H PD_H[3] PD_H[2] PD_H[1] PD_H[0]
+ PDEN_H_N[1] PDEN_H_N[0] PGHS_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PUEN_H[1]
+ PUEN_H[0] PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0]
+ SLOW_H SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
*.PININFO DRVHI_H:I DRVLO_H_N:I I2C_MODE_H_N:I NGHS_H:I OE_I_H_N:I
*.PININFO PAD:B PD_DIS_H:I PD_H[3]:O PD_H[2]:O PD_H[1]:O PD_H[0]:O
*.PININFO PDEN_H_N[1]:I PDEN_H_N[0]:I PGHS_H:I PU_H_N[3]:O PU_H_N[2]:O
*.PININFO PU_H_N[1]:O PU_H_N[0]:O PUEN_H[1]:I PUEN_H[0]:I PUG_H:I
*.PININFO SLEW_CTL_H[1]:I SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I
*.PININFO SLEW_CTL_H_N[0]:I SLOW_H:I SLOW_H_N:I VCC_IO:I VGND_IO:I
*.PININFO VPB_DRVR:I VSSD:I
XI192 DRVLO_H_N en_cmos_b I2C_MODE_H_N NGHS_H nsw_en OE_I_H_N PAD PD_DIS_H
+ PD_H[3] PD_H[2] PDEN_H_N[1] PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0]
+ SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
+ sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix
XI191 DRVHI_H DRVLO_H_N en_cmos_b nsw_en PD_H[3] PD_H[2] PD_H[1] PD_H[0]
+ PDEN_H_N[1] PDEN_H_N[0] PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PUEN_H[1]
+ PUEN_H[0] SLOW_H SLOW_H_N VCC_IO VGND_IO sky130_fd_io__gpio_ovtv2_obpredrvr_old
.ENDS sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix DRVLO_H_N EN_CMOS_B
+ I2C_MODE_H_N NGHS_H NSW_EN OE_I_H_N PAD PD_DIS_H PD_H[3] PD_H[2] PDEN_H_N[1]
+ PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0]
+ SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
*.PININFO DRVLO_H_N:I EN_CMOS_B:O I2C_MODE_H_N:I NGHS_H:I NSW_EN:O
*.PININFO OE_I_H_N:I PAD:B PD_DIS_H:I PD_H[3]:O PD_H[2]:O
*.PININFO PDEN_H_N[1]:I PGHS_H:I PUG_H:I SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I
*.PININFO SLOW_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I VSSD:I
Xpd_strong_q0 DRVLO_H_N EN_CMOS_B I2C_MODE_H_N NGHS_H NSW_EN OE_I_H_N PAD
+ PD_DIS_H PD_H[3] PD_H[2] PDEN_H_N[1] PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0]
+ SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix
.ENDS sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_old DRVHI_H DRVLO_H_N EN_CMOS_B
+ NSW_EN PD_H[3] PD_H[2] PD_H[1] PD_H[0] PDEN_H_N[1] PDEN_H_N[0] PU_H_N[3]
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] PUEN_H[1] PUEN_H[0] SLOW_H SLOW_H_N VCC_IO VGND_IO
*.PININFO DRVHI_H:I DRVLO_H_N:I EN_CMOS_B:I NSW_EN:I PD_H[3]:O
*.PININFO PD_H[2]:O PD_H[1]:O PD_H[0]:O PDEN_H_N[1]:I PDEN_H_N[0]:I
*.PININFO PU_H_N[3]:O PU_H_N[2]:O PU_H_N[1]:O PU_H_N[0]:O PUEN_H[1]:I
*.PININFO PUEN_H[0]:I SLOW_H:I SLOW_H_N:I VCC_IO:I VGND_IO:I
xI19 VGND_IO VCC_IO sky130_fd_io__condiode
Xpu_strong_slow_q0 DRVHI_H PU_H_N[1] PUEN_H[1] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpu_weak_q0 DRVHI_H PU_H_N[0] PUEN_H[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_weak
XI151 DRVLO_H_N PD_H[0] PDEN_H_N[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_weak
Xpd_strong_slow_q0 DRVLO_H_N PD_H[1] EN_CMOS_B VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_strong_slow
XI150 DRVLO_H_N DRVLO_H_N EN_CMOS_B NSW_EN PD_H[3] PD_H[2] PDEN_H_N[1] SLOW_H
+ VCC_IO VGND_IO sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos
Xpu_strong_q0 DRVHI_H PU_H_N[3] PU_H_N[2] PUEN_H[1] SLOW_H_N VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong
.ENDS sky130_fd_io__gpio_ovtv2_obpredrvr_old

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix DM_H[2] DM_H[1]
+ DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] DRVHI_H HLD_I_H_N HLD_I_OVR_H NGHS_H
+ OD_I_H_N OE_HS_H OE_N OUT PAD PD_H[3] PD_H[2] PD_H[1] PD_H[0] PGHS_H PU_H_N[3]
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1]
+ SLEW_CTL_H_N[0] SLOW SLOW_H_N VCCD VDDIO VPB_DRVR VPWR_KA VSSD VSSIO
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I DRVHI_H:O HLD_I_H_N:I HLD_I_OVR_H:I NGHS_H:I
*.PININFO OD_I_H_N:I OE_HS_H:O OE_N:I OUT:I PAD:B PD_H[3]:O PD_H[2]:O
*.PININFO PD_H[1]:O PD_H[0]:O PGHS_H:I PU_H_N[3]:O PU_H_N[2]:O
*.PININFO PU_H_N[1]:O PU_H_N[0]:O PUG_H:I SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I SLOW:I
*.PININFO SLOW_H_N:O VCCD:I VDDIO:I VPB_DRVR:I VPWR_KA:I VSSD:I
*.PININFO VSSIO:I
Xpredrvr_q0 DRVHI_H drvlo_h_n pden_h_n<2> NGHS_H oe_i_h_n PAD net72 PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] pden_h_n<1> pden_h_n<0> PGHS_H PU_H_N[3] PU_H_N[2]
+ PU_H_N[1] PU_H_N[0] puen_h<1> puen_h<0> PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0]
+ SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] slow_h SLOW_H_N VDDIO VSSIO VPB_DRVR VSSD
+ sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix
Xdatoe_q0 DRVHI_H drvlo_h_n HLD_I_H_N HLD_I_OVR_H OD_I_H_N oe_h OE_N OUT net72
+ VDDIO VSSD VPWR_KA sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix
Xctl_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N OD_I_H_N
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> net86 net85 puen_h<1> puen_h<0> SLOW slow_h
+ SLOW_H_N VDDIO VSSD VCCD VDDIO sky130_fd_io__gpio_ovtv2_octl_i2c_fix
XI354 oe_hs_i_h oe_hs_i_h_n VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x1
XI353 oe_h oe_i_h_n VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x2
XI355 oe_hs_i_h_n OE_HS_H VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x2
XI351 net86 net85 n<1> VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_nor
XI352 n<1> oe_i_h_n oe_hs_i_h VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_nor
.ENDS sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_octl_i2c_fix DM_H[2] DM_H[1] DM_H[0] DM_H_N[2]
+ DM_H_N[1] DM_H_N[0] HLD_I_H_N OD_I_H_N PDEN_H_N[2] PDEN_H_N[1] PDEN_H_N[0]
+ PUEN_0_H PUEN_2OR1_H PUEN_H[1] PUEN_H[0] SLOW SLOW_H SLOW_H_N VCC_IO VGND VPWR
+ VREG_EN_H_N
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I OD_I_H_N:I PDEN_H_N[2]:O
*.PININFO PDEN_H_N[1]:O PDEN_H_N[0]:O PUEN_0_H:O PUEN_2OR1_H:O
*.PININFO PUEN_H[1]:O PUEN_H[0]:O SLOW:I SLOW_H:O SLOW_H_N:O VCC_IO:I
*.PININFO VGND:I VPWR:I VREG_EN_H_N:I
XI211 n<8> DM_H_N[1] PUEN_0_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI201 DM_H_N[2] DM_H_N[1] n<9> VGND VCC_IO sky130_fd_io__hvsbt_nor
XI366 DM_H[1] DM_H[0] net87 VGND VCC_IO sky130_fd_io__hvsbt_nor
XI210 DM_H[2] DM_H[0] n<8> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI200 DM_H[2] DM_H[1] n<10> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI185 DM_H_N[0] n<4> net207 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI186 DM_H_N[2] DM_H_N[1] n<4> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI187 DM_H[1] DM_H[0] n<3> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI208 PUEN_2OR1_H VREG_EN_H_N n<5> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI203 n<10> DM_H[0] n<1> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI204 n<9> DM_H_N[0] n<0> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> PUEN_2OR1_H VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI365 net87 DM_H[2] PDEN_H_N[2] VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n PUEN_H[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n PUEN_H[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 PDEN_H_N[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 PDEN_H_N[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI377 PUEN_0_H puen_h0_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI374 net207 pden_h1 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI381 OD_I_H_N n9 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xls_slow_q0 HLD_I_H_N SLOW SLOW_H SLOW_H_N n9 VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpio_ovtv2_octl_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix FORCE_H[1]
+ NGA_PAD_VPMP_H NGB_PAD_VPMP_H NGHS_H OD_I_H_N OE_HS_H PAD PD_CSD_H PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] PGHS_H PU_CSD_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0]
+ PUG_H[7] PUG_H[6] PUG_H[5] TIE_HI_ESD TIE_LO_ESD VDDIO VDDIO_AMX VPB_DRVR VSSA
+ VSSD VSSIO VSSIO_AMX
*.PININFO FORCE_H[1]:I NGA_PAD_VPMP_H:I NGB_PAD_VPMP_H:I NGHS_H:O
*.PININFO OD_I_H_N:I OE_HS_H:I PAD:O PD_CSD_H:I PD_H[3]:I PD_H[2]:I
*.PININFO PD_H[1]:I PD_H[0]:I PGHS_H:O PU_CSD_H:I PU_H_N[3]:I
*.PININFO PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I PUG_H[7]:B PUG_H[6]:B
*.PININFO PUG_H[5]:B TIE_HI_ESD:O TIE_LO_ESD:O VDDIO:I VDDIO_AMX:B
*.PININFO VPB_DRVR:B VSSA:I VSSD:I VSSIO:I VSSIO_AMX:I
Xhotswap_q0 FORCE_H[1] NGHS_H OD_I_H_N OE_HS_H p2g PAD pad_esd PGHS_H PUG_H[7]
+ PUG_H[6] PUG_H[5] pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> net74 VDDIO
+ VPB_DRVR VDDIO VSSD sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix
Xbondpad_q0 PAD VSSIO sky130_fd_io__com_pad
Xodrvr_q0 TIE_HI_ESD PAD pad_esd PD_CSD_H PD_H[3] PD_H[2] PD_H[1] PD_H[0] PGHS_H
+ PU_CSD_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] pug_h<4> pug_h<3> pug_h<2>
+ pug_h<1> pug_h<0> TIE_HI_ESD TIE_LO_ESD VDDIO VDDIO_AMX VPB_DRVR VSSD VSSIO
+ VSSIO_AMX sky130_fd_io__gpio_ovtv2_odrvr_sub
XI122<2> PD_H[3] PGHS_H net106<0> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI122<1> PD_H[2] PGHS_H net106<1> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI122<0> PD_H[1] PGHS_H net106<2> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85<2> net106<0> PGHS_H VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85<1> net106<1> PGHS_H VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85<0> net106<2> PGHS_H VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104<2> net102<0> PGHS_H VSSA VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104<1> net102<1> PGHS_H VSSA VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104<0> net102<2> PGHS_H VSSA VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI103<2> PD_CSD_H PGHS_H net102<0> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI103<1> NGA_PAD_VPMP_H PGHS_H net102<1> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI103<0> NGB_PAD_VPMP_H PGHS_H net102<2> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_sub NGHS_H PAD PAD_ESD PD_CSD_H PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] PGHS_H PU_CSD_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0]
+ PUG_H[4] PUG_H[3] PUG_H[2] PUG_H[1] PUG_H[0] TIE_HI_ESD TIE_LO_ESD VDDIO
+ VDDIO_AMX VPB_DRVR VSSD VSSIO VSSIO_AMX
*.PININFO NGHS_H:I PAD:B PAD_ESD:B PD_CSD_H:I PD_H[3]:I PD_H[2]:I
*.PININFO PD_H[1]:I PD_H[0]:I PGHS_H:I PU_CSD_H:I PU_H_N[3]:I
*.PININFO PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I PUG_H[4]:B PUG_H[3]:B
*.PININFO PUG_H[2]:B PUG_H[1]:B PUG_H[0]:B TIE_HI_ESD:B TIE_LO_ESD:B
*.PININFO VDDIO:I VDDIO_AMX:B VPB_DRVR:B VSSD:I VSSIO:I VSSIO_AMX:I
Xpddrvr_strong_slow_q0 strong_slow_pad PD_H[1] VDDIO VSSIO
+ sky130_fd_io__gpio_pddrvr_strong_slow
XI73 weak_pad PD_H[0] VDDIO VSSIO sky130_fd_io__gpio_pddrvr_weak
Xres_q0 strong_slow_pad PAD_ESD VSSIO sky130_fd_io__com_res_strong_slow
Xres_weak_q0 weak_pad PAD_ESD VSSIO sky130_fd_io__com_res_weak
Xpd_drvr_q0 PAD PD_CSD_H PD_H[3] PD_H[2] TIE_LO_ESD VDDIO VSSIO VSSIO_AMX
+ sky130_fd_io__gpio_ovtv2_pddrvr
Xpudrvr_weak_q0 NGHS_H weak_pad PGHS_H PU_H_N[0] PUG_H[0] VDDIO VPB_DRVR VSSD
+ VSSIO sky130_fd_io__gpio_ovtv2_pudrvr_weak
Xstrong_slow_pudrvr_q0 NGHS_H strong_slow_pad PGHS_H PU_H_N[1] PUG_H[1] VDDIO
+ VPB_DRVR VSSD VSSIO sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow
Xpudrvr_strong_q0 NGHS_H NGHS_H NGHS_H PAD PGHS_H PGHS_H PGHS_H PU_CSD_H
+ PU_H_N[3] PU_H_N[2] PUG_H[4] PUG_H[3] PUG_H[2] TIE_HI_ESD VDDIO VDDIO_AMX
+ VPB_DRVR VSSD VSSIO sky130_fd_io__gpio_ovtv2_pudrvr_strong
Xres_esd_q0 PAD_ESD PAD sky130_fd_io__res75only_small
xI72 VSSIO VDDIO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpio_ovtv2_odrvr_sub

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix DRVHI_H DRVLO_H_N HLD_H_N
+ HLD_I_OVR_H OD_I_H_N OE_H OE_N OUT PD_DIS_H VCC_IO VGND VPWR_KA
*.PININFO DRVHI_H:O DRVLO_H_N:O HLD_H_N:I HLD_I_OVR_H:I OD_I_H_N:I
*.PININFO OE_H:O OE_N:I OUT:I PD_DIS_H:O VCC_IO:I VGND:I VPWR_KA:I
Xdat_ls_q0 HLD_I_OVR_H OUT PD_DIS_H pu_dis_h VGND net60 VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls
Xcclat_q0 DRVHI_H DRVLO_H_N OE_H PD_DIS_H pu_dis_h VCC_IO VGND
+ sky130_fd_io__com_cclat_i2c_fix
XI36 OD_I_H_N net60 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI37 OD_I_H_N net56 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xoe_ls_q0 HLD_I_OVR_H OE_N OE_H net56 OD_I_H_N VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls_i2c_fix
.ENDS sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix DM_H[2] DM_H[1] DM_H[0]
+ DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N HLD_I_OVR_H NGA_PAD_VPMP_H
+ NGB_PAD_VPMP_H OD_I_H_N OE_N OUT PAD PD_CSD_H PGHS_H PU_CSD_H PUG_H[6] PUG_H[5]
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW TIE_HI_ESD
+ TIE_LO_ESD VCCD VDDIO VDDIO_AMX VPB_DRVR VPWR_KA VSSA VSSD VSSIO VSSIO_AMX
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I HLD_I_OVR_H:I NGA_PAD_VPMP_H:I
*.PININFO NGB_PAD_VPMP_H:I OD_I_H_N:I OE_N:I OUT:I PAD:O PD_CSD_H:I
*.PININFO PGHS_H:O PU_CSD_H:I PUG_H[6]:B PUG_H[5]:B SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I SLOW:I
*.PININFO TIE_HI_ESD:O TIE_LO_ESD:O VCCD:I VDDIO:I VDDIO_AMX:B
*.PININFO VPB_DRVR:B VPWR_KA:I VSSA:I VSSD:I VSSIO:I VSSIO_AMX:I
Xodrvr_q0 TIE_LO_ESD NGA_PAD_VPMP_H NGB_PAD_VPMP_H nghs_h OD_I_H_N oe_hs_h PAD
+ PD_CSD_H pd_h<3> pd_h<2> pd_h<1> pd_h<0> PGHS_H PU_CSD_H pu_h_n<3> pu_h_n<2>
+ pu_h_n<1> pu_h_n<0> pug_h<7> PUG_H[6] PUG_H[5] TIE_HI_ESD TIE_LO_ESD VDDIO
+ VDDIO_AMX VPB_DRVR VSSA VSSD VSSIO VSSIO_AMX
+ sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix
Xopath_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] drvhi_h
+ HLD_I_H_N HLD_I_OVR_H nghs_h OD_I_H_N oe_hs_h OE_N OUT PAD pd_h<3> pd_h<2>
+ pd_h<1> pd_h<0> PGHS_H pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<7>
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW slow_h_n VCCD
+ VDDIO VPB_DRVR VPWR_KA VSSD VSSIO
+ sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix
.ENDS sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr PAD PD_CSD PD_H[3] PD_H[2] TIE_LO_ESD
+ VDDIO VSSIO VSSIO_Q
*.PININFO PAD:B PD_CSD:I PD_H[3]:I PD_H[2]:I TIE_LO_ESD:O VDDIO:B
*.PININFO VSSIO:B VSSIO_Q:B
XI26 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xn1_q0 PAD PD_H[2] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn2_q0 PAD PD_H[2] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn3_q0 PAD PD_H[2] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn8_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn7_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn6_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn5_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn9_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn10_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn11_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
xI9 VSSIO VDDIO sky130_fd_io__condiode
xI62 VSSIO_Q VDDIO sky130_fd_io__condiode
* RI8 VDDIO net96 short	 ; This device does not exist. . .
Xn14_q0 PAD PD_CSD VSSIO_Q VSSIO_Q sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31
+ l=0.55 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xn13_q0 PAD PD_CSD VSSIO_Q VSSIO_Q sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31
+ l=0.55 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pddrvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr_unit ND NGIN NS
*.PININFO ND:B NGIN:I NS:B
Xndrv_q0 ND NGIN NS NS sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pddrvr_unit

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias DRVLO_H_N EN_H EN_H_N PBIAS
+ PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_H:I EN_H_N:I PBIAS:O PD_H:I PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
XE1 n<1> n<0> sky130_fd_io__tk_em1o
XE2 PBIAS pbias1 sky130_fd_io__tk_em1o
XE3 pbias1 net88 sky130_fd_io__tk_em1s
XE4 net108 PBIAS sky130_fd_io__tk_em1s
XE6 PBIAS net84 sky130_fd_io__tk_em1s
XE5 n<101> bias_g sky130_fd_io__tk_em1s
XI27 n<0> PD_H EN_H_N sky130_fd_io__tk_opto
XI47 PBIAS bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 n<1> DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 bias_g DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 n<0> n<0> n<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 drvlo_i_h DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 bias_g n<1> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 bias_g EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 net157 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 net108 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 n<1> PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI48 n<100> PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI41 n<101> PD_H n<100> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI44 PBIAS PBIAS pbias1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 pbias1 pbias1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net183 EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net171 n<0> net183 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 PBIAS EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 drvlo_i_h DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 bias_g DRVLO_H_N net171 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 PBIAS drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 N0 VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 net161 net161 N0 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net157 net157 net161 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net88 N0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI43 net84 bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI40 N0 drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos DRVHI_H DRVLO_H_N
+ EN_CMOS_B NSW_EN_INT PD_H[3] PD_H[2] PDEN_H_N SLOW_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I DRVLO_H_N:I EN_CMOS_B:I NSW_EN_INT:I PD_H[3]:O
*.PININFO PD_H[2]:O PDEN_H_N:I SLOW_H:I VCC_IO:I VGND_IO:I
Xbias_q0 DRVHI_H en_fast_h en_fast_h_n pbias_out PD_H[2] PDEN_H_N VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias
Xnr3_q0 DRVLO_H_N net76 net76 PD_H[2] NSW_EN_INT VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2
Xnr2_q0 DRVLO_H_N en_fast2_n<1> en_fast2_n<0> PD_H[3] NSW_EN_INT VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI76 net76 pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> VCC_IO sky130_fd_io__tk_opti
Xinv_q0 en_fast_h en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xnor_q0 SLOW_H EN_CMOS_B en_fast_h VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  Added 3rd terminal to res_generic_nd__hv devices

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix DRVLO_H_N EN_CMOS_B
+ I2C_MODE_H_N NGHS_H NSW_EN_INT OE_I_H_N PAD_CAP PD_DIS_H PD_H[3] PD_H[2]
+ PDEN_H_N[1] PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1]
+ SLEW_CTL_H_N[0] SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
*.PININFO DRVLO_H_N:I EN_CMOS_B:O I2C_MODE_H_N:I NGHS_H:I NSW_EN_INT:O
*.PININFO OE_I_H_N:I PAD_CAP:B PD_DIS_H:I PD_H[3]:O PD_H[2]:O
*.PININFO PDEN_H_N[1]:I PGHS_H:I PUG_H:I SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I
*.PININFO SLOW_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I VSSD:I
XI123 PD_DIS_H nsw_enb OE_I_H_N net200 VGND_IO VCC_IO sky130_fd_io__nor3_dnw
xI208 VGND_IO VCC_IO sky130_fd_io__condiode
XI161 net293 drvlo_h_n_i2c_2 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI159 net298 drvlo_h_n_i2c_1 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI224 net288 net247 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI605 en enb VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI176 net318 drvlo_h_n_i2c_4 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI191 nsw_en nsw_enb VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI198 net303 drvlo_h_n_i2c VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI179 net283 NSW_EN_INT VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI168 net263 mode1b VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI122 drvlo_h drvlo_h_n_buf VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI170 net278 mode3b VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI715 PDEN_H_N[1] pden_h<1> VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI162 net313 drvlo_h_n_i2c_3 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI254 DRVLO_H_N drvlo_h VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI602 vdelay net200 en VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
XI112 pden_h<1> nsw_enb EN_CMOS_B VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
XI430 SLEW_CTL_H[1] SLEW_CTL_H_N[0] net263 VGND_IO VCC_IO
+ sky130_fd_io__com_nand2_dnw
XI175 drvlo_h_n_i2c mode4b net318 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI163 drvlo_h_n_i2c mode3b net313 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI109 SLOW_H_N I2C_MODE_H_N nsw_en VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI197 nsw_enb drvlo_h_n_buf net303 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI158 drvlo_h_n_i2c mode1b net298 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI160 drvlo_h_n_i2c mode2b net293 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI225 SLEW_CTL_H[1] SLEW_CTL_H[0] net288 VGND_IO VCC_IO
+ sky130_fd_io__com_nor2_dnw
XI181 PDEN_H_N[1] nsw_en net283 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI169 SLEW_CTL_H[1] SLEW_CTL_H_N[0] net278 VGND_IO VCC_IO
+ sky130_fd_io__com_nor2_dnw
XI94 nsw_en nsw_enb PD_H[2] PD_H[3] VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_predrvr_switch
XI288 N0 net193 VSSD sky130_fd_pr__res_generic_nd__hv W=0.5 L=113.375 m=1
XI287 vdiode net190 VSSD sky130_fd_pr__res_generic_nd__hv W=0.5 L=113.375 m=1
XI206 N0 en VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI190 net531 en VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI220 net420 enb VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI153 PD_H[2] PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI182 VGND_IO vdelay VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0
+ l=2.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI201 net352 N0 net190 VGND_IO sky130_fd_pr__nfet_05v0_nvt m=10 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI625 net404 PD_H[3] net348 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI339 net400 pden_h<1> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI125 PD_H[3] drvlo_h_n_buf net400 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI344 PD_H[3] PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI63 net388 vdiode PD_H[3] VGND_IO sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI189 net388 VGND_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI10 biasp vdiode net336 VGND_IO sky130_fd_pr__nfet_05v0_nvt m=5 w=10.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI374 net519 nsw_en PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI137 biasp1 vdiode VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 net369 net369 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 vdiode vdiode VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI165 vdiode en VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 N0 N0 net369 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net352 N0 net190 VGND_IO sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI755 net348 PD_H[3] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI579 vdelay drvlo_h net404 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI192 net519 VGND_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI219 net336 vdiode vr VGND_IO sky130_fd_pr__nfet_01v8_lvt m=5 w=7.0 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI232<1> cas3 PGHS_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI232<0> cas10 PGHS_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI278 VGND_IO VGND_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 PUG_H NGHS_H nsw_enb VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI245 cas10 VCC_IO cas4 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI196 nc biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=5 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI200 cas3 biasp1 nc VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI199 PD_H[3] drvlo_h_n_i2c_2 cas3 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI205 net352 en VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI156 cas5 biasp1 ne VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI580 vdelay drvlo_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI136 biasp biasp1 na VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI144 cas4 biasp1 nd VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI84 PD_H[3] drvlo_h_n_i2c cas2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI230 nc VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI79 nb biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=17 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI260 net535 enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI228 PD_H[3] drvlo_h_n_i2c net535 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI73 net388 drvlo_h_n_i2c net531 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI561 PD_H[3] drvlo_h_n_i2c_1 cas4 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI560 nd biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=14 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI375 PD_H[3] PUG_H net519 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI164 biasp enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI167 biasp1 enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI138 biasp1 biasp1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI145 cas2 biasp1 nb VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI141 na biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=10 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI154 ne biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=14 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI178 net193 en VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI155 PD_H[3] drvlo_h_n_i2c_3 cas5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI241 cas10 biasp1 nf VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI240 nf biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=8 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI229 ne VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=4.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI217 nb VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=3 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI216 nd VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI215 cas3 VCC_IO cas2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI214 cas5 VCC_IO cas2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI239 PD_H[3] drvlo_h_n_i2c_3 cas10 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI213 cas3 VCC_IO cas4 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI212 na VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI211 VCC_IO VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=4 w=0.55 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI210 VCC_IO VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=6 w=0.55 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<5> na enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<4> nb enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<3> nc enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<2> nd enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<1> ne enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<0> nf enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 nsw_enb PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI70 net531 en VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XRI221 net420 vr sky130_fd_pr__res_generic_po W=0.75 L=513.445 m=1
RI186 SLEW_CTL_H_N[0] mode4b sky130_fd_pr__res_generic_m1 L=0.035 W=1
RI157 net247 mode2b sky130_fd_pr__res_generic_m1 L=0.035 W=1
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I PD_H:O PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xmnin_q0 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_slow_q0 PD_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_H DRVLO_H_N int_nor<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_H DRVLO_H_N int_nor<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast<1>_q0 int_nor<1> EN_FAST_N[1] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_fast<0>_q0 int_nor<0> EN_FAST_N[0] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I PD_H:O PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xmnin_q0 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_slow_q0 PD_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_H DRVLO_H_N int_nor<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_H DRVLO_H_N int_nor<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast<1>_q0 int_nor<1> EN_FAST_N[1] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_fast<0>_q0 int_nor<0> EN_FAST_N[0] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_predrvr_switch NMOS_EN PMOS_EN SIG1 SIG2 VCC_IO
+ VGND_IO
*.PININFO NMOS_EN:I PMOS_EN:I SIG1:B SIG2:B VCC_IO:I VGND_IO:I
XI374 SIG1 NMOS_EN SIG2 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI375 SIG2 PMOS_EN SIG1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_predrvr_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong NGHS_H[4] NGHS_H[3] NGHS_H[2] PAD
+ PGHS_H[4] PGHS_H[3] PGHS_H[2] PU_CSD_H PU_H_N[3] PU_H_N[2] PUG_H[4] PUG_H[3]
+ PUG_H[2] TIE_HI_ESD VDDIO VDDIO_AMX VPB_DRVR VSSD VSSIO
*.PININFO NGHS_H[4]:I NGHS_H[3]:I NGHS_H[2]:I PAD:B PGHS_H[4]:I
*.PININFO PGHS_H[3]:I PGHS_H[2]:I PU_CSD_H:I PU_H_N[3]:I PU_H_N[2]:I
*.PININFO PUG_H[4]:B PUG_H[3]:B PUG_H[2]:B TIE_HI_ESD:O VDDIO:I
*.PININFO VDDIO_AMX:B VPB_DRVR:B VSSD:I VSSIO:I
XI49 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
XI133 VPB_DRVR tie_hi_vpbdrvr sky130_fd_io__tk_tie_r_out_esd
XI112 PUG_H[2] net83 sky130_fd_io__tk_em2o
XI111 PUG_H[4] net81 sky130_fd_io__tk_em1o
XI141 PUG_H[3] net79 sky130_fd_io__tk_em2o
XI152 PUG_H[4] net079 sky130_fd_io__tk_em2o
XI142 tie_hi_vpbdrvr net79 sky130_fd_io__tk_em2s
XI82 tie_hi_vpbdrvr net83 sky130_fd_io__tk_em2s
XI109 tie_hi_vpbdrvr net81 sky130_fd_io__tk_em2s
XI153 tie_hi_vpbdrvr net079 sky130_fd_io__tk_em2s
Xn7_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn6_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<2>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<1>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<0>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn4_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<3>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<2>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<1>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<0>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<1>_q0 VPB_DRVR PAD net79 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<0>_q0 VPB_DRVR PAD net79 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<1>_q0 VPB_DRVR PAD PUG_H[4] VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<0>_q0 VPB_DRVR PAD PUG_H[4] VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<1>_q0 VPB_DRVR PAD net81 VDDIO_AMX sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<0>_q0 VPB_DRVR PAD net81 VDDIO_AMX sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<1>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<0>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<1>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<0>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<1>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<0>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<1>_q0 VPB_DRVR PAD net079 VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<0>_q0 VPB_DRVR PAD net079 VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
XI136 PUG_H[4] NGHS_H[4] PU_CSD_H VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI127 PUG_H[2] NGHS_H[2] PU_H_N[2] VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 PUG_H[3] NGHS_H[3] PU_H_N[3] VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI137 PU_CSD_H PGHS_H[4] PUG_H[4] VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI128 PU_H_N[2] PGHS_H[2] PUG_H[2] VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI24 PU_H_N[3] PGHS_H[3] PUG_H[3] VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow NGHS_H PAD PGHS_H PU_H_N
+ PUG_H VDDIO VPB_DRVR VSSD VSSIO
*.PININFO NGHS_H:I PAD:B PGHS_H:I PU_H_N:I PUG_H:B VDDIO:I VPB_DRVR:I
*.PININFO VSSD:I VSSIO:I
XI20 PUG_H NGHS_H PU_H_N VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 PU_H_N PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpdrv_q0 PAD PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=12 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5 PB PD PGIN PS
*.PININFO PB:B PD:B PGIN:I PS:B
Xpdrv_q0 PD PGIN PS PB sky130_fd_pr__esd_pfet_g5v0d10v5 m=1 w=15.5 l=0.55 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_weak NGHS_H PAD PGHS_H PU_H_N PUG_H
+ VDDIO VPB_DRVR VSSD VSSIO
*.PININFO NGHS_H:I PAD:B PGHS_H:I PU_H_N:I PUG_H:B VDDIO:I VPB_DRVR:I
*.PININFO VSSD:I VSSIO:I
XI36 PAD net26 sky130_fd_io__tk_em2o
XI51 PUG_H NGHS_H PU_H_N VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI50 PU_H_N PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpdrv_q0 PAD PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=3 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 net26 PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 PAD PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong DRVHI_H PU_H_N[3] PU_H_N[2]
+ PUEN_H SLOW_H_N VCC_IO VGND_IO
*.PININFO DRVHI_H:I PU_H_N[3]:O PU_H_N[2]:O PUEN_H:I SLOW_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xnd2b_q0 DRVHI_H en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0>
+ PU_H_N[3] PUEN_H VCC_IO VGND_IO sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3
Xnd2a_q0 DRVHI_H net54 net54 net54 net54 PU_H_N[2] PUEN_H VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h sky130_fd_io__tk_opto
Xinv_q0 en_fast_h_n en_fast_h VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xnbias_q0 DRVHI_H en_fast_h en_fast_h_n nbias_out PU_H_N[2] PUEN_H VCC_IO
+ VGND_IO sky130_fd_io__com_pupredrvr_nbias
Xnand_q0 PUEN_H SLOW_H_N en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
.ENDS sky130_fd_io__gpio_ovtv2_pupredrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2 DRVHI_H EN_FAST[3]
+ EN_FAST[2] EN_FAST[1] EN_FAST[0] PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_FAST[3]:I EN_FAST[2]:I EN_FAST[1]:I
*.PININFO EN_FAST[0]:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XE1 net30 PU_H_N sky130_fd_io__tk_em1s
XRrespu1 int_res net30 sky130_fd_pr__res_generic_po W=0.33 L=11 m=1
XRrespu2 PU_H_N int_res sky130_fd_pr__res_generic_po W=0.33 L=4 m=1
Xmnin_fast<3>_q0 net30 DRVHI_H int<3> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<2>_q0 net30 DRVHI_H int<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<1>_q0 net30 DRVHI_H int<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<0>_q0 net30 DRVHI_H int<0> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_slow1_q0 n<2> PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.75 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_slow_q0 PU_H_N DRVHI_H n<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_fast<3>_q0 int<3> EN_FAST[3] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<2>_q0 int<2> EN_FAST[2] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<1>_q0 int<1> EN_FAST[1] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<0>_q0 int<0> EN_FAST[0] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_q0 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_q0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3 DRVHI_H EN_FAST[3]
+ EN_FAST[2] EN_FAST[1] EN_FAST[0] PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_FAST[3]:I EN_FAST[2]:I EN_FAST[1]:I
*.PININFO EN_FAST[0]:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XE1 net30 PU_H_N sky130_fd_io__tk_em1s
XRrespu1 int_res net30 sky130_fd_pr__res_generic_po W=0.33 L=11 m=1
XRrespu2 PU_H_N int_res sky130_fd_pr__res_generic_po W=0.33 L=4 m=1
Xmnin_fast<3>_q0 net30 DRVHI_H int<3> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<2>_q0 net30 DRVHI_H int<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<1>_q0 net30 DRVHI_H int<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<0>_q0 net30 DRVHI_H int<0> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_slow1_q0 n<2> PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.75 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_slow_q0 PU_H_N DRVHI_H n<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_fast<3>_q0 int<3> EN_FAST[3] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<2>_q0 int<2> EN_FAST[2] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<1>_q0 int<1> EN_FAST[1] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<0>_q0 int<0> EN_FAST[0] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_q0 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_q0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pddrvr_strong FORCE_LO_H FORCE_LOVOL_H PAD PD_H[3]
+ PD_H[2] TIE_LO_ESD VCC_IO VGND_IO VSSIO_AMX
*.PININFO FORCE_LO_H:I FORCE_LOVOL_H:I PAD:O PD_H[3]:I PD_H[2]:I
*.PININFO TIE_LO_ESD:O VCC_IO:I VGND_IO:I VSSIO_AMX:I
XI112 PD_H[2] net61 sky130_fd_io__tk_em2s
XI113 PD_H[2] net59 sky130_fd_io__tk_em2s
XI97 PD_H[3] net85 sky130_fd_io__tk_em2s
XI108 TIE_LO_ESD net83 sky130_fd_io__tk_em2s
XI109 TIE_LO_ESD net77 sky130_fd_io__tk_em2s
XI102 PD_H[3] net73 sky130_fd_io__tk_em2s
XI104 PD_H[3] net69 sky130_fd_io__tk_em2s
XI96 PD_H[3] net67 sky130_fd_io__tk_em2s
XI87 TIE_LO_ESD net59 sky130_fd_io__tk_em2o
XI83 PD_H[3] net61 sky130_fd_io__tk_em2o
XI99 TIE_LO_ESD net85 sky130_fd_io__tk_em2o
XI82 TIE_LO_ESD net61 sky130_fd_io__tk_em2o
XI98 PD_H[2] net85 sky130_fd_io__tk_em2o
XI106 PD_H[2] net83 sky130_fd_io__tk_em2o
XI107 PD_H[3] net83 sky130_fd_io__tk_em2o
XI110 PD_H[3] net77 sky130_fd_io__tk_em2o
XI111 PD_H[2] net77 sky130_fd_io__tk_em2o
XI100 TIE_LO_ESD net73 sky130_fd_io__tk_em2o
XI101 PD_H[2] net73 sky130_fd_io__tk_em2o
XI103 TIE_LO_ESD net69 sky130_fd_io__tk_em2o
XI105 PD_H[2] net69 sky130_fd_io__tk_em2o
XI95 PD_H[2] net67 sky130_fd_io__tk_em2o
XI94 TIE_LO_ESD net67 sky130_fd_io__tk_em2o
XI88 PD_H[3] net59 sky130_fd_io__tk_em2o
XI49 VGND_IO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xn24<2>_q0 PAD net85 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1>_q0 PAD net85 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0>_q0 PAD net85 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2>_q0 PAD net67 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1>_q0 PAD net67 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0>_q0 PAD net67 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn12_q0 PAD net61 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2>_q0 PAD net69 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1>_q0 PAD net69 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0>_q0 PAD net69 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2>_q0 PAD net83 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1>_q0 PAD net83 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0>_q0 PAD net83 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn13_q0 PAD net59 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn31_q0 PAD net73 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
xI72 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpio_pddrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pddrvr_strong_slow PAD PD_H VCC_IO VGND_IO
*.PININFO PAD:O PD_H:I VCC_IO:I VGND_IO:I
Xndrv_q0 PAD PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_pddrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pddrvr_weak PAD PD_H VCC_IO VGND_IO
*.PININFO PAD:O PD_H:I VCC_IO:I VGND_IO:I
Xndrv1_q0 PAD PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_pddrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pudrvr_strong PAD PU_H_N[3] PU_H_N[2] TIE_HI_ESD
+ VCC_IO VNB
*.PININFO PAD:O PU_H_N[3]:I PU_H_N[2]:I TIE_HI_ESD:O VCC_IO:I VNB:I
XI112 PU_H_N[2] net43 sky130_fd_io__tk_em2s
XI108 TIE_HI_ESD net59 sky130_fd_io__tk_em2s
XI109 TIE_HI_ESD net53 sky130_fd_io__tk_em2s
XI104 PU_H_N[3] net49 sky130_fd_io__tk_em2s
XI125 PU_H_N[3] net45 sky130_fd_io__tk_em2s
XI83 PU_H_N[3] net43 sky130_fd_io__tk_em2o
XI82 TIE_HI_ESD net43 sky130_fd_io__tk_em2o
XI106 PU_H_N[2] net59 sky130_fd_io__tk_em2o
XI107 PU_H_N[3] net59 sky130_fd_io__tk_em2o
XI110 PU_H_N[3] net53 sky130_fd_io__tk_em2o
XI111 PU_H_N[2] net53 sky130_fd_io__tk_em2o
XI103 TIE_HI_ESD net49 sky130_fd_io__tk_em2o
XI105 PU_H_N[2] net49 sky130_fd_io__tk_em2o
XI124 TIE_HI_ESD net45 sky130_fd_io__tk_em2o
XI123 PU_H_N[2] net45 sky130_fd_io__tk_em2o
XI49 VCC_IO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xn24<2>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<1>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<0>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<2>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<1>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<0>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn22_q0 PAD net45 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn21_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<2>_q0 PAD net43 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<1>_q0 PAD net43 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<0>_q0 PAD net43 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<2>_q0 PAD net49 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<1>_q0 PAD net49 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<0>_q0 PAD net49 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<1>_q0 PAD net59 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<0>_q0 PAD net59 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<2>_q0 PAD net53 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<1>_q0 PAD net53 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<0>_q0 PAD net53 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<2>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<1>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<0>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<2>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<1>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<0>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<2>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<1>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<0>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
.ENDS sky130_fd_io__gpio_pudrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pudrvr_unit_2_5 PD PGIN PS
*.PININFO PD:B PGIN:I PS:B
Xpdrv_q0 PD PGIN PS PS sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_pudrvr_unit_2_5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL
+ ANALOG_SEL ENABLE_VDDA_H ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N OUT PAD VCCD VDDA
+ VDDIO_Q VSSA VSSD VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I ENABLE_VDDA_H:I ENABLE_VSWITCH_H:I HLD_I_H:I
*.PININFO HLD_I_H_N:I OUT:I PAD:B VCCD:I VDDA:I VDDIO_Q:I VSSA:I
*.PININFO VSSD:I VSSIO_Q:I VSWITCH:I
xI43 VSSIO_Q VDDA sky130_fd_io__condiode
xI78 VSSA VSWITCH sky130_fd_io__condiode
Xmux_a_q0 AMUXBUS_A nga_amx_vpmp_h nga_pad_vpmp_h nmida_vccd net101 net101 net97
+ net97 net100 net99 net0127 HLD_I_H pga_amx_vdda_h_n pga_pad_vddioq_h_n VDDA
+ VDDIO_Q VSSA VSSD sky130_fd_io__gpiov2_amux_switch
Xmux_b_q0 AMUXBUS_B ngb_amx_vpmp_h ngb_pad_vpmp_h nmidb_vccd net101 net101 net97
+ net97 net100 net99 net0127 HLD_I_H pgb_amx_vdda_h_n pgb_pad_vddioq_h_n VDDA
+ VDDIO_Q VSSA VSSD sky130_fd_io__gpiov2_amux_switch
XBBM_logic ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H net0127
+ ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N nga_amx_vpmp_h nga_pad_vpmp_h ngb_amx_vpmp_h
+ ngb_pad_vpmp_h nmida_vccd nmidb_vccd OUT pd_csd_vswitch_h pga_amx_vdda_h_n
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n VCCD
+ VDDA VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_ctl_logic
XI26 PAD net99 sky130_fd_io__res75only_small
XI58 net168 net97 sky130_fd_io__res75only_small
XI28 net166 net101 sky130_fd_io__res75only_small
XI57 PAD net168 sky130_fd_io__res75only_small
XI27 PAD net100 sky130_fd_io__res75only_small
XI55 PAD PAD sky130_fd_io__res75only_small
XI54 PAD net166 sky130_fd_io__res75only_small
XI53 PAD PAD sky130_fd_io__res75only_small
XI39 PAD net81 sky130_fd_io__res75only_small
XI40 PAD net85 sky130_fd_io__res75only_small
XI52 net81 pu_csd_vddioq_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=3
+ w=15.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XMP_PU net85 pu_csd_vddioq_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=4
+ w=15.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI49 net81 pd_csd_vswitch_h VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 m=6
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XMN_PD net85 pd_csd_vswitch_h VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 m=8
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI27 OUT IN VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 OUT IN VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_inv_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic ANALOG_EN ANALOG_POL ANALOG_SEL
+ ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N
+ NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H
+ NMIDA_VCCD NMIDB_VCCD OUT PD_CSD_VSWITCH_H PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N VCCD VDDA VDDIO_Q VSSA
+ VSSD VSWITCH
*.PININFO ANALOG_EN:I ANALOG_POL:I ANALOG_SEL:I ENABLE_VDDA_H:I
*.PININFO ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I HLD_I_H:I HLD_I_H_N:I
*.PININFO NGA_AMX_VSWITCH_H:O NGA_PAD_VSWITCH_H:O NGB_AMX_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H:O NMIDA_VCCD:O NMIDB_VCCD:O OUT:I
*.PININFO PD_CSD_VSWITCH_H:O PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O
*.PININFO PGB_AMX_VDDA_H_N:O PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
Xamux_sw_drvr_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h
+ amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on
+ amuxbusa_on_n amuxbusb_on amuxbusb_on_n NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H
+ nga_pad_vswitch_h_n NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n
+ nmida_on_n NMIDA_VCCD nmida_vccd_n nmidb_on_n NMIDB_VCCD nmidb_vccd_n
+ PD_CSD_VSWITCH_H pd_csd_vswitch_h_n pd_on pd_on_n PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N pu_on
+ pu_on_n VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_drvr
Xamux_lv_decoder_q0 amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n
+ ANALOG_EN ANALOG_POL ANALOG_SEL NGA_PAD_VSWITCH_H nga_pad_vswitch_h_n
+ NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n
+ nmidb_vccd_n OUT pd_on pd_on_n pd_csd_vswitch_h_n PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N pu_on pu_on_n
+ PU_CSD_VDDIOQ_H_N VCCD VSSD sky130_fd_io__gpiov2_amux_decoder
Xamux_ls_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n
+ amux_en_vswitch_h amux_en_vswitch_h_n ANALOG_EN ENABLE_VDDA_H ENABLE_VDDA_H_N
+ ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
+ sky130_fd_io__gpiov2_amux_ls
.ENDS sky130_fd_io__gpiov2_amux_ctl_logic

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix ANALOG_EN ANALOG_POL
+ ANALOG_SEL ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H_N
+ NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H
+ NMIDA_VCCD NMIDB_VCCD OUT PD_CSD_VSWITCH_H PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N VCCD VDDA VDDIO_Q VSSA
+ VSSD VSWITCH
*.PININFO ANALOG_EN:I ANALOG_POL:I ANALOG_SEL:I ENABLE_VDDA_H:I
*.PININFO ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I HLD_I_H_N:I
*.PININFO NGA_AMX_VSWITCH_H:O NGA_PAD_VSWITCH_H:O NGB_AMX_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H:O NMIDA_VCCD:O NMIDB_VCCD:O OUT:I
*.PININFO PD_CSD_VSWITCH_H:O PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O
*.PININFO PGB_AMX_VDDA_H_N:O PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
Xamux_ls_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vswitch_h
+ amux_en_vswitch_h_n ANALOG_EN ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H
+ HLD_I_H_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
+ sky130_fd_io__gpiov2_amux_ls_i2c_fix
Xamux_sw_drvr_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h
+ amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on amuxbusa_on_n amuxbusb_on
+ amuxbusb_on_n HLD_I_H_N NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H nga_pad_vswitch_h_n
+ NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n nmida_on_n NMIDA_VCCD
+ nmida_vccd_n nmidb_on_n NMIDB_VCCD nmidb_vccd_n PD_CSD_VSWITCH_H
+ pd_csd_vswitch_h_n pd_on pd_on_n PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N pu_on pu_on_n VCCD VDDA
+ VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_drvr_i2c_fix
Xamux_lv_decoder_q0 amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n
+ ANALOG_EN ANALOG_POL ANALOG_SEL NGA_PAD_VSWITCH_H nga_pad_vswitch_h_n
+ NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n
+ nmidb_vccd_n OUT pd_on pd_on_n pd_csd_vswitch_h_n PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N pu_on pu_on_n
+ PU_CSD_VDDIOQ_H_N VCCD VSSD sky130_fd_io__gpiov2_amux_decoder
.ENDS sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls IN IN_B OUT_H OUT_H_N RST_H RST_H_N
+ VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST_H:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I VPWR_LV:I
XI14 OUT_H fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H_N fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 net61 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI58 fbk VPWR_LV net62 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI59 fbk_n VPWR_LV net66 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net66 IN net61 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net62 IN_B net61 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix IN IN_B OUT_H RST_H RST_H_N
+ VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O RST_H:I RST_H_N:I VGND:I VPWR_HV:I
*.PININFO VPWR_LV:I
XI14 fbk_n RST_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 net70 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI58 fbk VPWR_LV net71 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI59 fbk_n VPWR_LV net75 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net75 IN net70 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net71 IN_B net70 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_lshv2hv IN IN_B OUT_H OUT_H_N RST_H
+ RST_H_N VGND VPWR_HV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST_H:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I
XI14 OUT_H_N fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI64 net64 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 fbk_n IN net64 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 fbk IN_B net64 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_lshv2hv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_decoder AMUXBUSA_ON AMUXBUSA_ON_N AMUXBUSB_ON
+ AMUXBUSB_ON_N ANALOG_EN ANALOG_POL ANALOG_SEL NGA_PAD_VSWITCH_H
+ NGA_PAD_VSWITCH_H_N NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N NMIDA_ON_N
+ NMIDA_VCCD_N D_B NMIDB_VCCD_N OUT PD_ON PD_ON_N PD_VSWITCH_H_N PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_ON PU_ON_N
+ PU_VDDIOQ_H_N VCCD VSSD
*.PININFO AMUXBUSA_ON:O AMUXBUSA_ON_N:O AMUXBUSB_ON:O AMUXBUSB_ON_N:O
*.PININFO ANALOG_EN:I ANALOG_POL:I ANALOG_SEL:I NGA_PAD_VSWITCH_H:I
*.PININFO NGA_PAD_VSWITCH_H_N:I NGB_PAD_VSWITCH_H:I
*.PININFO NGB_PAD_VSWITCH_H_N:I NMIDA_ON_N:O NMIDA_VCCD_N:I D_B:O
*.PININFO NMIDB_VCCD_N:I OUT:I PD_ON:O PD_ON_N:O PD_VSWITCH_H_N:I
*.PININFO PGA_AMX_VDDA_H_N:I PGA_PAD_VDDIOQ_H_N:I PGB_AMX_VDDA_H_N:I
*.PININFO PGB_PAD_VDDIOQ_H_N:I PU_ON:O PU_ON_N:O PU_VDDIOQ_H_N:I
*.PININFO VCCD:I VSSD:I
XI116 ana_en_i_n int_pd_on_n int_pd_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI113 ana_en_i_n net144 int_amuxa_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI115 ana_en_i_n int_pu_on_n int_pu_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI114 ana_en_i_n net137 int_amuxb_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI111 ana_pol_i out_i int_pu_on_n VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI112 ana_pol_i_n out_i_n int_pd_on_n VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI109 ana_sel_i_n pol_xor_out net144 VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI110 pol_xor_out ana_sel_i net137 VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI106 NGB_PAD_VSWITCH_H net212 net172 VSSD VCCD sky130_fd_io__hvsbt_nor
XI102 NGA_PAD_VSWITCH_H net222 net167 VSSD VCCD sky130_fd_io__hvsbt_nor
XI79 int_pu_on PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H_N
+ NGB_PAD_VSWITCH_H_N int_fbk_puon_n VSSD VCCD sky130_fd_io__gpiov2_amux_nand5
XI80 int_pd_on PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H_N
+ NGB_PAD_VSWITCH_H_N int_fbk_pdon_n VSSD VCCD sky130_fd_io__gpiov2_amux_nand5
XI78 int_amuxb_on PU_VDDIOQ_H_N PD_VSWITCH_H_N NMIDB_VCCD_N AMUXBUSB_ON_N VSSD
+ VCCD sky130_fd_io__gpiov2_amux_nand4
XI77 int_amuxa_on PU_VDDIOQ_H_N PD_VSWITCH_H_N NMIDA_VCCD_N AMUXBUSA_ON_N VSSD
+ VCCD sky130_fd_io__gpiov2_amux_nand4
XI101 PGA_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N net222 VSSD VCCD
+ sky130_fd_io__hvsbt_nand2
XI121 int_amux_b_on_n net172 D_B VSSD VCCD sky130_fd_io__hvsbt_nand2
XI105 PGB_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N net212 VSSD VCCD
+ sky130_fd_io__hvsbt_nand2
XI120 int_amux_a_on_n net167 NMIDA_ON_N VSSD VCCD sky130_fd_io__hvsbt_nand2
XI45 ana_pol_i out_i pol_xor_out VSSD VCCD sky130_fd_io__xor2_1
XI41 ana_pol_i_n ana_pol_i VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI89 int_amuxa_on int_amux_a_on_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI39 ANALOG_SEL ana_sel_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI40 ana_sel_i_n ana_sel_i VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI35 ANALOG_POL ana_pol_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI74 AMUXBUSB_ON_N AMUXBUSB_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI73 AMUXBUSA_ON_N AMUXBUSA_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI76 int_fbk_pdon_n PD_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI58 ANALOG_EN ana_en_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI75 int_fbk_puon_n PU_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI43 OUT out_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI44 out_i_n out_i VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI91 int_amuxb_on int_amux_b_on_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI93 PU_ON PU_ON_N VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI95 PD_ON PD_ON_N VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
.ENDS sky130_fd_io__gpiov2_amux_decoder

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N
+ AMUXBUSA_ON AMUXBUSA_ON_N AMUXBUSB_ON AMUXBUSB_ON_N NGA_AMX_VSWITCH_H
+ NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H
+ NGB_PAD_VSWITCH_H_N NMIDA_ON_N NMIDA_VCCD NMIDA_VCCD_N D_B NMIDB_VCCD
+ NMIDB_VCCD_N PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N PD_ON PD_ON_N PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N PU_ON
+ PU_ON_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:I AMUX_EN_VDDA_H_N:I AMUX_EN_VDDIO_H:I
*.PININFO AMUX_EN_VDDIO_H_N:I AMUX_EN_VSWITCH_H:I
*.PININFO AMUX_EN_VSWITCH_H_N:I AMUXBUSA_ON:I AMUXBUSA_ON_N:I
*.PININFO AMUXBUSB_ON:I AMUXBUSB_ON_N:I NGA_AMX_VSWITCH_H:O
*.PININFO NGA_PAD_VSWITCH_H:O NGA_PAD_VSWITCH_H_N:O
*.PININFO NGB_AMX_VSWITCH_H:O NGB_PAD_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H_N:O NMIDA_ON_N:I NMIDA_VCCD:O
*.PININFO NMIDA_VCCD_N:O D_B:I NMIDB_VCCD:O NMIDB_VCCD_N:O
*.PININFO PD_CSD_VSWITCH_H:O PD_CSD_VSWITCH_H_N:O PD_ON:I PD_ON_N:I
*.PININFO PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O PGB_AMX_VDDA_H_N:O
*.PININFO PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O PU_ON:I PU_ON_N:I
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
XI93 NMIDA_VCCD NMIDA_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
XI105 NMIDB_VCCD NMIDB_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
XI38 net274 PU_CSD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_pucsd_inv
Xpga_amx_ls_q0 net265 net272 PGA_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H
+ VSSA VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net239 net245 PGB_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H VSSA VDDA
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net256 NGA_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI42 net265 PGA_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI47 net256 NGA_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI62 net239 PGB_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI63 net236 NGB_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI64 net236 NGB_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI53 D_B NMIDB_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
XI89 NMIDA_ON_N NMIDA_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv_q0 net254 PD_CSD_VSWITCH_H VSWITCH VSSA
+ sky130_fd_io__gpiov2_amx_pdcsd_inv
XI90 PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI85 NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI87 NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
Xpu_csd_ls_q0 PU_ON PU_ON_N net274 net275 AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H VSSD
+ VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpga_pad_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net265 net272 AMUX_EN_VDDIO_H_N
+ AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xnga_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net257 net256 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls_q0 PD_ON PD_ON_N net248 net254 AMUX_EN_VSWITCH_H_N AMUX_EN_VSWITCH_H
+ VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpgb_pad_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net239 net245 AMUX_EN_VDDIO_H_N
+ AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net230 net236 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
XI76 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI77 NGB_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI75 NGA_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI78 NGA_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI104 PD_CSD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_i2c_fix AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N AMUXBUSA_ON AMUXBUSA_ON_N
+ AMUXBUSB_ON AMUXBUSB_ON_N HLD_I_H_N NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H
+ NGA_PAD_VSWITCH_H_N NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N
+ NMIDA_ON_N NMIDA_VCCD NMIDA_VCCD_N D_B NMIDB_VCCD NMIDB_VCCD_N PD_CSD_VSWITCH_H
+ PD_CSD_VSWITCH_H_N PD_ON PD_ON_N PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N PU_ON PU_ON_N VCCD VDDA
+ VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:I AMUX_EN_VDDA_H_N:I AMUX_EN_VDDIO_H:I
*.PININFO AMUX_EN_VSWITCH_H:I AMUX_EN_VSWITCH_H_N:I AMUXBUSA_ON:I
*.PININFO AMUXBUSA_ON_N:I AMUXBUSB_ON:I AMUXBUSB_ON_N:I HLD_I_H_N:I
*.PININFO NGA_AMX_VSWITCH_H:O NGA_PAD_VSWITCH_H:O
*.PININFO NGA_PAD_VSWITCH_H_N:O NGB_AMX_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H:O NGB_PAD_VSWITCH_H_N:O NMIDA_ON_N:I
*.PININFO NMIDA_VCCD:O NMIDA_VCCD_N:O D_B:I NMIDB_VCCD:O
*.PININFO NMIDB_VCCD_N:O PD_CSD_VSWITCH_H:O PD_CSD_VSWITCH_H_N:O
*.PININFO PD_ON:I PD_ON_N:I PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O
*.PININFO PGB_AMX_VDDA_H_N:O PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O
*.PININFO PU_ON:I PU_ON_N:I VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I
*.PININFO VSWITCH:I
Xpga_pad_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net154 net160 hld_i_h HLD_I_H_N
+ amux_en_vddio_h_n AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
Xpgb_pad_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net144 net149 hld_i_h HLD_I_H_N
+ amux_en_vddio_h_n AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
XI38 net168 PU_CSD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_pucsd_buf
Xpu_csd_ls_q0 PU_ON PU_ON_N net167 net168 HLD_I_H_N AMUX_EN_VDDIO_H VSSD VDDIO_Q
+ VCCD sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3
XI111 HLD_I_H_N hld_i_h VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI110 AMUX_EN_VDDIO_H amux_en_vddio_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI93 NMIDA_VCCD NMIDA_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
XI105 NMIDB_VCCD NMIDB_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
Xpga_amx_ls_q0 net154 net160 PGA_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H
+ VSSA VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net144 net149 PGB_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H VSSA VDDA
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net295 NGA_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI42 net154 PGA_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI47 net295 NGA_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI62 net144 PGB_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI63 net284 NGB_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI64 net284 NGB_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI53 D_B NMIDB_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
XI89 NMIDA_ON_N NMIDA_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv_q0 net293 PD_CSD_VSWITCH_H VSWITCH VSSA
+ sky130_fd_io__gpiov2_amx_pdcsd_inv
XI87 NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI85 NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI90 PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
Xnga_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net296 net295 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls_q0 PD_ON PD_ON_N net287 net293 AMUX_EN_VSWITCH_H_N AMUX_EN_VSWITCH_H
+ VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net278 net284 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
XI76 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI77 NGB_PAD_VSWITCH_H amux_en_vddio_h_n VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI75 NGA_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI78 NGA_PAD_VSWITCH_H amux_en_vddio_h_n VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI104 PD_CSD_VSWITCH_H amux_en_vddio_h_n VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls IN IN_B OUT_H OUT_H_N RST_H RST_H_N
+ VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST_H:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I VPWR_LV:I
XI11 OUT_H_N OUT_H VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 net42 VPWR_LV net58 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 net38 VPWR_LV net54 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net58 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net54 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT_H RST_H_N net38 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 OUT_H_N RST_H_N net42 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3 IN IN_B OUT_H OUT_H_N
+ RST2_H_N RST_H_N VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST2_H_N:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I VPWR_LV:I
XI34 RST_H_N net086 VGND VPWR_HV sky130_fd_io__hvsbt_inv_x1
XI33 RST2_H_N net074 VGND VPWR_HV sky130_fd_io__hvsbt_inv_x1
XI11 OUT_H_N OUT_H VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 OUT_H_N RST2_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 OUT_H_N RST_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 net55 VPWR_LV net79 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 net51 VPWR_LV net75 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 OUT_H net086 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net79 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net75 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 OUT_H net074 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT_H RST_H_N net51 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 OUT_H_N RST_H_N net55 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2 IN IN_B OUT_H OUT_H_N
+ RST2_H RST2_H_N RST_H RST_H_N VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST2_H:I RST2_H_N:I RST_H:I
*.PININFO RST_H_N:I VGND:I VPWR_HV:I VPWR_LV:I
XI11 OUT_H_N OUT_H VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 OUT_H_N RST2_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 OUT_H_N RST_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 net56 VPWR_LV net76 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 net52 VPWR_LV net72 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net76 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net72 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 OUT_H RST2_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT_H RST_H_N net52 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 OUT_H_N RST_H_N net56 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_lshv2hv IN IN_B OUT_H_N RST_H RST_H_N
+ VGND VPWR_HV
*.PININFO IN:I IN_B:I OUT_H_N:O RST_H:I RST_H_N:I VGND:I VPWR_HV:I
XI14 OUT_H_N fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI64 net52 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 fbk_n IN net52 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 fbk IN_B net52 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_lshv2hv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ls AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N
+ ANALOG_EN ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N VCCD
+ VDDA VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:O AMUX_EN_VDDA_H_N:O AMUX_EN_VDDIO_H:O
*.PININFO AMUX_EN_VDDIO_H_N:O AMUX_EN_VSWITCH_H:O
*.PININFO AMUX_EN_VSWITCH_H_N:O ANALOG_EN:I ENABLE_VDDA_H:I
*.PININFO ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I HLD_I_H:I HLD_I_H_N:I
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
XI32 ENABLE_VDDA_H ENABLE_VDDA_H_N VSSA VDDA sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls_q0 AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VSWITCH_H
+ AMUX_EN_VSWITCH_H_N net74 ENABLE_VSWITCH_H VSSA VSWITCH
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls_q0 AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ ENABLE_VDDA_H_N ENABLE_VDDA_H VSSA VDDA sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 ANALOG_EN ana_en_i_n VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 ENABLE_VSWITCH_H net74 VSSA VSWITCH sky130_fd_io__hvsbt_inv_x1
Xpd_vddio_ls_q0 ana_en_i ana_en_i_n AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N HLD_I_H
+ HLD_I_H_N VSSD VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_ctl_ls
.ENDS sky130_fd_io__gpiov2_amux_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ls_i2c_fix AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N ANALOG_EN ENABLE_VDDA_H
+ ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:O AMUX_EN_VDDA_H_N:O AMUX_EN_VDDIO_H:O
*.PININFO AMUX_EN_VSWITCH_H:O AMUX_EN_VSWITCH_H_N:O ANALOG_EN:I
*.PININFO ENABLE_VDDA_H:I ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I
*.PININFO HLD_I_H_N:I VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
Xpd_vddio_ls_q0 ana_en_i ana_en_i_n AMUX_EN_VDDIO_H net082 HLD_I_H_N VSSD
+ VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix
XI32 ENABLE_VDDA_H ENABLE_VDDA_H_N VSSA VDDA sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls_q0 AMUX_EN_VDDIO_H net028 AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N
+ net83 ENABLE_VSWITCH_H VSSA VSWITCH sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls_q0 AMUX_EN_VDDIO_H net028 AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ ENABLE_VDDA_H_N ENABLE_VDDA_H VSSA VDDA sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 ANALOG_EN ana_en_i_n VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 ENABLE_VSWITCH_H net83 VSSA VSWITCH sky130_fd_io__hvsbt_inv_x1
XI36 AMUX_EN_VDDIO_H net028 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI35 HLD_I_H_N net082 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_amux_ls_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ls_inv_x1 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ls_inv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_nand4 IN0 IN1 IN2 IN3 OUT VGND VPWR
*.PININFO IN0:I IN1:I IN2:I IN3:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 out_n OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 OUT out_n VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net50 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net58 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net54 IN3 net58 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 net50 IN2 net54 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 out_n OUT VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 VGND out_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_nand4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_nand5 IN0 IN1 IN2 IN3 IN4 OUT VGND VPWR
*.PININFO IN0:I IN1:I IN2:I IN3:I IN4:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 OUT out_n VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 out_n OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net51 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 net63 IN4 net59 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net59 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net55 IN3 net63 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 net51 IN2 net55 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 out_n OUT VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 VGND out_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_nand5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_switch AMUXBUS_HV NG_AMX_VPMP_H NG_PAD_VPMP_H
+ NMID_VCCD PAD_HV_N0 PAD_HV_N1 PAD_HV_N2 PAD_HV_N3 PAD_HV_P0 PAD_HV_P1 PD_H_VDDA
+ PD_H_VDDIO PG_AMX_VDDA_H_N PG_PAD_VDDIOQ_H_N VDDA VDDIO VSSA VSSD
*.PININFO AMUXBUS_HV:B NG_AMX_VPMP_H:I NG_PAD_VPMP_H:I NMID_VCCD:I
*.PININFO PAD_HV_N0:B PAD_HV_N1:B PAD_HV_N2:B PAD_HV_N3:B PAD_HV_P0:B
*.PININFO PAD_HV_P1:B PD_H_VDDA:I PD_H_VDDIO:I PG_AMX_VDDA_H_N:I
*.PININFO PG_PAD_VDDIOQ_H_N:I VDDA:I VDDIO:I VSSA:I VSSD:I
xI72 VSSA VDDA sky130_fd_io__condiode
xI71 mid1 VDDA sky130_fd_io__condiode
xI70 mid VDDA sky130_fd_io__condiode
XI56 VSSA net79 sky130_fd_io__res75only_small
XI12 VSSA net77 sky130_fd_io__res75only_small
XI46 PAD_HV_N3 NG_PAD_VPMP_H mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 mid NG_PAD_VPMP_H PAD_HV_N1 mid sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 PAD_HV_N0 NG_PAD_VPMP_H mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 mid1 NG_PAD_VPMP_H PAD_HV_N2 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 mid NG_AMX_VPMP_H AMUXBUS_HV mid sky130_fd_pr__nfet_g5v0d10v5 m=7 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI57 mid1 NMID_VCCD net79 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI47 mid1 NG_AMX_VPMP_H AMUXBUS_HV mid1 sky130_fd_pr__nfet_g5v0d10v5 m=7 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI78<1> mid PD_H_VDDA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI78<0> mid1 PD_H_VDDA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77<1> mid PD_H_VDDIO VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77<0> mid1 PD_H_VDDIO VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 mid NMID_VCCD net77 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 mid PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 m=5 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 mid PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=3
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI36 mid PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=3
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_inv4 A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI75 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_inv4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_pdcsd_inv A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI414 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI519 Y VSSA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI517 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.0 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI429 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.0 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_pdcsd_inv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_buf A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI75 int A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.42 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 Y int VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=3 w=0.42 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74 int A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 Y int VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=5 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_pucsd_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_inv A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI75 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=7 w=0.42 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=7 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_pucsd_inv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ctl DM[2] DM[1] DM[0] DM_H[2] DM_H[1] DM_H[0]
+ DM_H_N[2] DM_H_N[1] DM_H_N[0] ENABLE_H ENABLE_INP_H HLD_H_N HLD_I_H HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS
+ INP_DIS_H_N OD_I_H VCC_IO VGND VPWR VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O ENABLE_H:I
*.PININFO ENABLE_INP_H:I HLD_H_N:I HLD_I_H:O HLD_I_H_N:O HLD_I_OVR_H:O
*.PININFO HLD_OVR:I IB_MODE_SEL:I IB_MODE_SEL_H:O IB_MODE_SEL_H_N:O
*.PININFO INP_DIS:I INP_DIS_H_N:O OD_I_H:O VCC_IO:I VGND:I VPWR:I
*.PININFO VTRIP_SEL:I VTRIP_SEL_H:O VTRIP_SEL_H_N:O
XI75 ENABLE_INP_H ENABLE_H startup_rst_h VGND VCC_IO sky130_fd_io__hvsbt_nor
Xhld_dis_blk_q0 ENABLE_H HLD_H_N HLD_I_H HLD_I_H_N HLD_I_OVR_H HLD_OVR OD_I_H
+ VCC_IO VGND VPWR sky130_fd_io__gpiov2_ctl_hld
Xls_bank_q0 DM[2] DM[1] DM[0] DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS net80
+ INP_DIS_H_N OD_I_H startup_rst_h inp_startup_en_h VCC_IO VGND VPWR VTRIP_SEL
+ VTRIP_SEL_H VTRIP_SEL_H_N sky130_fd_io__gpiov2_ctl_lsbank
XI56 OD_I_H ENABLE_INP_H net92 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI57 net92 inp_startup_en_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_ctl

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ctl_hld ENABLE_H HLD_H_N HLD_I_H HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR OD_I_H VCC_IO VGND VPWR
*.PININFO ENABLE_H:I HLD_H_N:I HLD_I_H:O HLD_I_H_N:O HLD_I_OVR_H:O
*.PININFO HLD_OVR:I OD_I_H:O VCC_IO:I VGND:I VPWR:I
Xhld_ovr_ls_q0 net65 HLD_OVR hld_ovr_h net37 od_h VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
XI30 OD_I_H hld_i_ovr_h_n HLD_I_OVR_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI26 net65 hld_ovr_h hld_i_ovr_h_n VGND VCC_IO sky130_fd_io__hvsbt_nor
Xhld_i_h_inv4_q0 net65 enable_vdda_h_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x4
XI31 od_i_h_n OD_I_H VGND VCC_IO sky130_fd_io__hvsbt_inv_x4
Xhld_nand_q0 ENABLE_H HLD_H_N net64 VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xod_h_inv_q0 ENABLE_H od_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv1_q0 net64 net65 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI32 od_h od_i_h_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv8<1>_q0 enable_vdda_h_n hld_i_h_n_net<1> VGND VCC_IO
+ sky130_fd_io__hvsbt_inv_x8
Xhld_i_h_inv8<0>_q0 enable_vdda_h_n hld_i_h_n_net<0> VGND VCC_IO
+ sky130_fd_io__hvsbt_inv_x8
* Rshort<1> hld_i_h_n_net<1> HLD_I_H_N short
* Rshort<0> hld_i_h_n_net<0> HLD_I_H_N short
* Rshort_hld_i_h enable_vdda_h_n HLD_I_H short
Rshort<1> hld_i_h_n_net<1> HLD_I_H_N sky130_fd_pr__res_generic_m1 L=1 W=1
Rshort<0> hld_i_h_n_net<0> HLD_I_H_N sky130_fd_pr__res_generic_m1 L=1 W=1
Rshort_hld_i_h enable_vdda_h_n HLD_I_H sky130_fd_pr__res_generic_m1 L=1 W=1
.ENDS sky130_fd_io__gpiov2_ctl_hld

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ctl_lsbank DM[2] DM[1] DM[0] DM_H[2] DM_H[1]
+ DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N IB_MODE_SEL IB_MODE_SEL_H
+ IB_MODE_SEL_H_N INP_DIS INP_DIS_H INP_DIS_H_N OD_I_H STARTUP_RST_H STARTUP_ST_H
+ VCC_IO VGND VPWR VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O HLD_I_H_N:I
*.PININFO IB_MODE_SEL:I IB_MODE_SEL_H:O IB_MODE_SEL_H_N:O INP_DIS:I
*.PININFO INP_DIS_H:O INP_DIS_H_N:O OD_I_H:I STARTUP_RST_H:I
*.PININFO STARTUP_ST_H:I VCC_IO:I VGND:I VPWR:I VTRIP_SEL:I
*.PININFO VTRIP_SEL_H:O VTRIP_SEL_H_N:O
Xtrip_sel_st_q0 trip_sel_st_h OD_I_H VGND sky130_fd_io__tk_opti
Xtrip_sel_rst_q0 trip_sel_rst_h VGND OD_I_H sky130_fd_io__tk_opti
Xie_n_rst_q0 ie_n_rst_h STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_opti
Xie_n_st_q0 ie_n_st_h STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> OD_I_H VGND sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> OD_I_H VGND sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> VGND OD_I_H sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> VGND OD_I_H sky130_fd_io__tk_opti
* NOTE:  This has the selectable open and short on metal2 instead of metal1
XI598 ib_mode_sel_st_h OD_I_H VGND sky130_fd_io__tk_optiB
* NOTE:  This has the selectable short on metal2 instead of metal1
XI597 ib_mode_sel_rst_h VGND OD_I_H sky130_fd_io__tk_optiA
XI337<1> dm_st_h<0> STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_opti
Xdm_ls<0>_q0 HLD_I_H_N DM[0] DM_H[0] DM_H_N[0] dm_rst_h<0> dm_st_h<0> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
Xinp_dis_ls_q0 HLD_I_H_N INP_DIS INP_DIS_H INP_DIS_H_N ie_n_rst_h ie_n_st_h
+ VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xtrip_sel_ls_q0 HLD_I_H_N VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N trip_sel_rst_h
+ trip_sel_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<2>_q0 HLD_I_H_N DM[2] DM_H[2] DM_H_N[2] dm_rst_h<2> dm_st_h<2> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<1>_q0 HLD_I_H_N DM[1] DM_H[1] DM_H_N[1] dm_rst_h<1> dm_st_h<1> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
XI595 HLD_I_H_N IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N ib_mode_sel_rst_h
+ ib_mode_sel_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpiov2_ctl_lsbank

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ibuf_se ENABLE_VDDIO_LV IBUFMUX_OUT IBUFMUX_OUT_H
+ IN_H IN_VT MODE_NORMAL_N MODE_VCCHIB_N VCCHIB VDDIO_Q VSSD VTRIP_SEL_H
+ VTRIP_SEL_H_N
*.PININFO ENABLE_VDDIO_LV:I IBUFMUX_OUT:O IBUFMUX_OUT_H:O IN_H:I
*.PININFO IN_VT:I MODE_NORMAL_N:I MODE_VCCHIB_N:I VCCHIB:I VDDIO_Q:I
*.PININFO VSSD:I VTRIP_SEL_H:I VTRIP_SEL_H_N:I
XI148 ENABLE_VDDIO_LV mode_vcchib mode_vcchib_lv_n VSSD VCCHIB
+ sky130_fd_io__hvsbt_nand2
XI149 ENABLE_VDDIO_LV mode_normal mode_normal_lv_n VSSD VCCHIB
+ sky130_fd_io__hvsbt_nand2
XI112 mode_normal_lv_n mode_normal_lv VSSD VSSD VCCHIB VCCHIB
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1
XI111 mode_vcchib_lv_n mode_vcchib_lv VSSD VSSD VCCHIB VCCHIB
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xlvls_q0 out_vcchib out_vddio mode_normal_lv mode_normal_lv_n mode_vcchib_lv
+ mode_vcchib_lv_n IBUFMUX_OUT net57 VCCHIB VSSD sky130_fd_io__gpiov2_ipath_lvls
Xhvls_q0 out_vcchib out_vddio out_n_vcchib mode_normal MODE_NORMAL_N mode_vcchib
+ MODE_VCCHIB_N IBUFMUX_OUT_H net68 VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_hvls
XI88 IN_H mode_vcchib_lv_n out_vcchib out_n_vcchib VCCHIB VSSD
+ sky130_fd_io__gpiov2_vcchib_in_buf
Xbuf_q0 IN_H IN_VT MODE_NORMAL_N out_vddio out_n_vddio VDDIO_Q VSSD VTRIP_SEL_H
+ VTRIP_SEL_H_N sky130_fd_io__gpiov2_in_buf
XI491 MODE_NORMAL_N mode_normal VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI105 MODE_VCCHIB_N mode_vcchib VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_ibuf_se

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ictl_logic DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS_H_N INP_DIS_I_H INP_DIS_I_H_N
+ MODE_NORMAL_N MODE_VCCHIB_N TRIPSEL_I_H TRIPSEL_I_H_N VDDIO_Q VSSD VTRIP_SEL_H_N
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I IB_MODE_SEL_H:I
*.PININFO IB_MODE_SEL_H_N:I INP_DIS_H_N:I INP_DIS_I_H:O
*.PININFO INP_DIS_I_H_N:O MODE_NORMAL_N:O MODE_VCCHIB_N:O
*.PININFO TRIPSEL_I_H:O TRIPSEL_I_H_N:O VDDIO_Q:I VSSD:I
*.PININFO VTRIP_SEL_H_N:I
XI71 VTRIP_SEL_H_N MODE_NORMAL_N TRIPSEL_I_H VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
XI80 dm_buf_dis_n INP_DIS_H_N INP_DIS_I_H VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI79 DM_H_N[2] and_dm01 dm_buf_dis_n VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI78 DM_H_N[1] DM_H_N[0] nand_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI36 INP_DIS_I_H_N IB_MODE_SEL_H MODE_VCCHIB_N VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
XI35 INP_DIS_I_H_N IB_MODE_SEL_H_N MODE_NORMAL_N VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
XI111 INP_DIS_I_H INP_DIS_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI75 nand_dm01 and_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI74 TRIPSEL_I_H TRIPSEL_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_ictl_logic

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_in_buf IN_H IN_VT MODE_NORMAL_N OUT OUT_N VDDIO_Q
+ VSSD VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO IN_H:I IN_VT:I MODE_NORMAL_N:I OUT:O OUT_N:O VDDIO_Q:I
*.PININFO VSSD:I VTRIP_SEL_H:I VTRIP_SEL_H_N:I
XI43 mode_normal_cmos_h mode_normal_cmos_h_n VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_inv_x1
XI488 VTRIP_SEL_H MODE_NORMAL_N mode_normal_cmos_h VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
XI583 IN_VT VTRIP_SEL_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI644 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI646 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI593 net91 MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI592 net103 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI591 fbk IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI590 fbk2 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI589 net91 in_b VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI588 fbk IN_VT VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI587 in_b IN_H fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI586 OUT_N net91 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI642 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI629 in_b IN_H net158 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI636 net158 mode_normal_cmos_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI632 net122 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI647 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.8 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI600 net103 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI598 net91 in_b net138 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI597 fbk2 mode_normal_cmos_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI596 OUT_N net91 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI595 net138 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI631 in_b IN_H net122 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI643 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_inbuf_lvinv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ipath DM_H_N[2] DM_H_N[1] DM_H_N[0] ENABLE_VDDIO_LV
+ IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS_H_N OUT OUT_H PAD VCCHIB VDDIO_Q VSSD
+ VTRIP_SEL_H_N
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I ENABLE_VDDIO_LV:I
*.PININFO IB_MODE_SEL_H:I IB_MODE_SEL_H_N:I INP_DIS_H_N:I OUT:O
*.PININFO OUT_H:O PAD:B VCCHIB:I VDDIO_Q:I VSSD:I VTRIP_SEL_H_N:I
XI106 ENABLE_VDDIO_LV OUT OUT_H in_h in_vt mode_normal_n mode_vcchib_n VCCHIB
+ VDDIO_Q VSSD tripsel_i_h tripsel_i_h_n sky130_fd_io__gpiov2_ibuf_se
XI107 DM_H_N[2] DM_H_N[1] DM_H_N[0] IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS_H_N
+ en_h_n en_h mode_normal_n mode_vcchib_n tripsel_i_h tripsel_i_h_n VDDIO_Q VSSD
+ VTRIP_SEL_H_N sky130_fd_io__gpiov2_ictl_logic
XI120 PAD in_h in_vt VDDIO_Q VSSD tripsel_i_h
+ sky130_fd_io__gpio_ovtv2_buf_localesd
.ENDS sky130_fd_io__gpiov2_ipath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ipath_hvls IN_VCCHIB IN_VDDIO INB_VCCHIB
+ MODE_NORMAL MODE_NORMAL_N MODE_VCCHIB MODE_VCCHIB_N OUT OUT_B VDDIO_Q VSSD
*.PININFO IN_VCCHIB:I IN_VDDIO:I INB_VCCHIB:I MODE_NORMAL:I
*.PININFO MODE_NORMAL_N:I MODE_VCCHIB:I MODE_VCCHIB_N:I OUT:O OUT_B:O
*.PININFO VDDIO_Q:I VSSD:I
XI325 fbk fbk_b VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI324 fbk_b fbk VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI323 net63 MODE_NORMAL VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI322 OUT_B IN_VDDIO net75 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI321 net75 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI320 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI319 OUT_B MODE_VCCHIB net63 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI318 net55 MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI317 OUT_B net84 net55 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI336 net84 fbk_b VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI335 OUT_B net84 net88 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI334 fbk INB_VCCHIB net116 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI333 net116 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI332 net112 MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI331 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI330 OUT_B IN_VDDIO net112 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI329 fbk_b IN_VCCHIB net92 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI328 fbk MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI327 net92 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI326 net88 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI337 net84 fbk_b VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_ipath_hvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ipath_lvls IN_VCCHIB IN_VDDIO MODE_NORMAL_LV
+ MODE_NORMAL_LV_N MODE_VCCHIB_LV MODE_VCCHIB_LV_N OUT OUT_B VCCHIB VSSD
*.PININFO IN_VCCHIB:I IN_VDDIO:I MODE_NORMAL_LV:I MODE_NORMAL_LV_N:I
*.PININFO MODE_VCCHIB_LV:I MODE_VCCHIB_LV_N:I OUT:O OUT_B:O VCCHIB:I
*.PININFO VSSD:I
XI345 fbk_n IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI344 net70 MODE_VCCHIB_LV VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI343 OUT_B fbk net78 VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI342 net78 MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI341 OUT_B MODE_NORMAL_LV net70 VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI340 net50 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI339 fbk_n MODE_NORMAL_LV VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI338 fbk fbk_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI337 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=4 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI336 OUT_B IN_VCCHIB net50 VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI351 net111 MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI350 OUT_B fbk net111 VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI349 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI348 fbk fbk_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI347 net95 MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI346 OUT_B IN_VCCHIB net95 VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI353 fbk_n IN_VDDIO net115 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI352 net115 MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_ipath_lvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_obpredrvr DRVHI_H DRVLO_H_N I2C_MODE_H_N PD_H[4]
+ PD_H[3] PD_H[2] PD_H[1] PD_H[0] PDEN_H_N[1] PDEN_H_N[0] PU_H_N[3] PU_H_N[2]
+ PU_H_N[1] PU_H_N[0] PUEN_H[1] PUEN_H[0] SLOW_H SLOW_H_N TIE_HI_ESD VCC_IO VGND
+ VGND_IO
*.PININFO DRVHI_H:I DRVLO_H_N:I I2C_MODE_H_N:I PD_H[4]:O PD_H[3]:O
*.PININFO PD_H[2]:O PD_H[1]:O PD_H[0]:O PDEN_H_N[1]:I PDEN_H_N[0]:I
*.PININFO PU_H_N[3]:O PU_H_N[2]:O PU_H_N[1]:O PU_H_N[0]:O PUEN_H[1]:I
*.PININFO PUEN_H[0]:I SLOW_H:I SLOW_H_N:I TIE_HI_ESD:I VCC_IO:I VGND:I
*.PININFO VGND_IO:I
Xpu_strong_q0 DRVHI_H PU_H_N[3] PU_H_N[2] PUEN_H[1] SLOW_H_N VCC_IO VGND_IO
+ sky130_fd_io__gpiov2_pupredrvr_strong
Xpd_strong_q0 DRVLO_H_N I2C_MODE_H_N PD_H[4] PD_H[3] PD_H[2] PDEN_H_N[1] SLOW_H
+ TIE_HI_ESD VCC_IO VGND VGND_IO sky130_fd_io__gpiov2_pdpredrvr_strong
Xpu_weak_q0 DRVHI_H PU_H_N[0] PUEN_H[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_weak
Xpd_weak_q0 DRVLO_H_N PD_H[0] PDEN_H_N[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_weak
Xpu_strong_slow_q0 DRVHI_H PU_H_N[1] PUEN_H[1] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpd_strong_slow_q0 DRVLO_H_N PD_H[1] PDEN_H_N[1] VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_strong_slow
xI15 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpiov2_obpredrvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_octl DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N OD_H PDEN_H_N[2] PDEN_H_N[1] PDEN_H_N[0] PUEN_0_H
+ PUEN_2OR1_H PUEN_H[1] PUEN_H[0] SLOW SLOW_H SLOW_H_N VCC_IO VGND VPWR
+ VREG_EN_H_N
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I OD_H:I PDEN_H_N[2]:O PDEN_H_N[1]:O
*.PININFO PDEN_H_N[0]:O PUEN_0_H:O PUEN_2OR1_H:O PUEN_H[1]:O
*.PININFO PUEN_H[0]:O SLOW:I SLOW_H:O SLOW_H_N:O VCC_IO:I VGND:I
*.PININFO VPWR:I VREG_EN_H_N:I
XI211 n<8> DM_H_N[1] PUEN_0_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI201 DM_H_N[2] DM_H_N[1] n<9> VGND VCC_IO sky130_fd_io__hvsbt_nor
XI381 DM_H[1] DM_H[0] net70 VGND VCC_IO sky130_fd_io__hvsbt_nor
XI210 DM_H[2] DM_H[0] n<8> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI200 DM_H[2] DM_H[1] n<10> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI185 DM_H_N[0] n<4> net130 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI186 DM_H_N[2] DM_H_N[1] n<4> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI187 DM_H[1] DM_H[0] n<3> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI208 PUEN_2OR1_H VREG_EN_H_N n<5> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI203 n<10> DM_H[0] n<1> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI204 n<9> DM_H_N[0] n<0> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> PUEN_2OR1_H VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI382 DM_H[2] net70 PDEN_H_N[2] VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n PUEN_H[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n PUEN_H[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 PDEN_H_N[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 PDEN_H_N[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI377 PUEN_0_H puen_h0_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI374 net130 pden_h1 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xls_slow_q0 HLD_I_H_N SLOW SLOW_H SLOW_H_N OD_H VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpiov2_octl

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_octl_dat DM_H[2] DM_H[1] DM_H[0] DM_H_N[2]
+ DM_H_N[1] DM_H_N[0] DRVHI_H HLD_I_H_N HLD_I_OVR_H OD_H OE_N OUT PD_H[4] PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] SLOW SLOW_H_N
+ TIE_HI_ESD VCC_IO VGND VGND_IO VPWR VPWR_KA
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I DRVHI_H:O HLD_I_H_N:I HLD_I_OVR_H:I OD_H:I
*.PININFO OE_N:I OUT:I PD_H[4]:O PD_H[3]:O PD_H[2]:O PD_H[1]:O
*.PININFO PD_H[0]:O PU_H_N[3]:O PU_H_N[2]:O PU_H_N[1]:O PU_H_N[0]:O
*.PININFO SLOW:I SLOW_H_N:O TIE_HI_ESD:I VCC_IO:I VGND:I VGND_IO:I
*.PININFO VPWR:I VPWR_KA:I
Xdatoe_q0 DRVHI_H drvlo_h_n HLD_I_H_N HLD_I_OVR_H OD_H oe_h OE_N OUT VCC_IO VGND
+ VPWR_KA sky130_fd_io__gpiov2_opath_datoe
Xctl_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N OD_H
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0>
+ SLOW slow_h SLOW_H_N VCC_IO VGND VPWR VCC_IO sky130_fd_io__gpiov2_octl
Xpredrvr_q0 DRVHI_H drvlo_h_n pden_h_n<2> PD_H[4] PD_H[3] PD_H[2] PD_H[1]
+ PD_H[0] pden_h_n<1> pden_h_n<0> PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0]
+ puen_h<1> puen_h<0> slow_h SLOW_H_N TIE_HI_ESD VCC_IO VGND VGND_IO
+ sky130_fd_io__gpiov2_obpredrvr
.ENDS sky130_fd_io__gpiov2_octl_dat

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_octl_mux A_H B_H SEL_H SEL_H_N VCCIO VSSIO Y_H
*.PININFO A_H:I B_H:I SEL_H:I SEL_H_N:I VCCIO:I VSSIO:I Y_H:O
XI2 Y_H SEL_H B_H VCCIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI3 Y_H SEL_H_N A_H VCCIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 B_H SEL_H_N Y_H VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 A_H SEL_H Y_H VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_octl_mux

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_odrvr FORCE_HI_H_N PAD PD_H[3] PD_H[2] PD_H[1]
+ PD_H[0] PD_H_I2C PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] TIE_HI_ESD TIE_LO_ESD
+ VCC_IO VGND VGND_IO
*.PININFO FORCE_HI_H_N:I PAD:O PD_H[3]:I PD_H[2]:I PD_H[1]:I PD_H[0]:I
*.PININFO PD_H_I2C:I PU_H_N[3]:I PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I
*.PININFO TIE_HI_ESD:O TIE_LO_ESD:O VCC_IO:I VGND:I VGND_IO:I
Xodrvr_q0 FORCE_HI_H_N PAD PD_H[3] PD_H[2] PD_H[1] PD_H[0] PD_H_I2C PU_H_N[3]
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] TIE_HI_ESD TIE_LO_ESD VCC_IO VGND VGND_IO
+ sky130_fd_io__gpiov2_odrvr_sub
Xbondpad_q0 PAD VGND_IO sky130_fd_io__com_pad
.ENDS sky130_fd_io__gpiov2_odrvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_odrvr_sub FORCE_HI_H_N PAD PD_H[3] PD_H[2] PD_H[1]
+ PD_H[0] PD_H_I2C PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] TIE_HI_ESD TIE_LO_ESD
+ VCC_IO VGND VGND_IO
*.PININFO FORCE_HI_H_N:I PAD:O PD_H[3]:I PD_H[2]:I PD_H[1]:I PD_H[0]:I
*.PININFO PD_H_I2C:I PU_H_N[3]:I PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I
*.PININFO TIE_HI_ESD:B TIE_LO_ESD:B VCC_IO:I VGND:I VGND_IO:I
Xpddrvr_strong_q0 PAD PD_H[3] PD_H[2] PD_H_I2C TIE_LO_ESD VCC_IO VGND_IO
+ sky130_fd_io__gpiov2_pddrvr_strong
Xpudrvr_strong_q0 PAD PU_H_N[3] PU_H_N[2] TIE_HI_ESD VCC_IO VGND
+ sky130_fd_io__gpio_pudrvr_strong
Xpudrvr_weak_q0 weak_pad PU_H_N[0] VCC_IO VGND VCC_IO
+ sky130_fd_io__com_pudrvr_weak
Xpddrvr_weak_q0 weak_pad PD_H[0] VCC_IO VGND_IO sky130_fd_io__gpio_pddrvr_weak
Xstrong_slow_pddrvr_q0 strong_slow_pad PD_H[1] VCC_IO VGND_IO
+ sky130_fd_io__gpio_pddrvr_strong_slow
Xstrong_slow_pudrvr_q0 strong_slow_pad PU_H_N[1] VCC_IO VGND VCC_IO
+ sky130_fd_io__com_pudrvr_strong_slow
Xres_q0 strong_slow_pad pad_r250 VGND_IO sky130_fd_io__com_res_strong_slow
Xres_weak_q0 weak_pad pad_r250 VGND_IO sky130_fd_io__com_res_weak
Xresd_q0 PAD pad_r250 sky130_fd_io__res250only_small
xI60 VGND_IO VCC_IO sky130_fd_io__condiode
xI59 VGND_IO VCC_IO sky130_fd_io__condiode
xI58 VGND_IO VCC_IO sky130_fd_io__condiode
xI72 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpiov2_odrvr_sub

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_opath DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N HLD_I_OVR_H OD_H OE_N OUT PAD SLOW TIE_HI_ESD TIE_LO_ESD
+ VCC_IO VGND VGND_IO VPWR VPWR_KA
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I HLD_I_OVR_H:I OD_H:I OE_N:I OUT:I
*.PININFO PAD:O SLOW:I TIE_HI_ESD:O TIE_LO_ESD:O VCC_IO:I VGND:I
*.PININFO VGND_IO:I VPWR:I VPWR_KA:I
Xodrvr_q0 net70 PAD pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h<4> pu_h_n<3> pu_h_n<2>
+ pu_h_n<1> pu_h_n<0> TIE_HI_ESD TIE_LO_ESD VCC_IO VGND VGND_IO
+ sky130_fd_io__gpiov2_odrvr
Xopath_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] drvhi_h
+ HLD_I_H_N HLD_I_OVR_H OD_H OE_N OUT pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0>
+ pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> SLOW slow_h_n TIE_HI_ESD VCC_IO VGND
+ VGND_IO VPWR VPWR_KA sky130_fd_io__gpiov2_octl_dat
.ENDS sky130_fd_io__gpiov2_opath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_opath_datoe DRVHI_H DRVLO_H_N HLD_H_N HLD_I_OVR_H
+ OD_H OE_H OE_N OUT VCC_IO VGND VPWR_KA
*.PININFO DRVHI_H:O DRVLO_H_N:O HLD_H_N:I HLD_I_OVR_H:I OD_H:I OE_H:O
*.PININFO OE_N:I OUT:I VCC_IO:I VGND:I VPWR_KA:I
Xdat_ls_q0 HLD_I_OVR_H OUT pd_dis_h pu_dis_h VGND OD_H VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls
Xoe_ls_q0 HLD_I_OVR_H OE_N oe_h_n OE_H VGND OD_H VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls
Xcclat_q0 DRVHI_H DRVLO_H_N oe_h_n pd_dis_h pu_dis_h VCC_IO VGND
+ sky130_fd_io__com_cclat
.ENDS sky130_fd_io__gpiov2_opath_datoe

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pddrvr_strong PAD PD_H[3] PD_H[2] PD_H_I2C
+ TIE_LO_ESD VCC_IO VGND_IO
*.PININFO PAD:O PD_H[3]:I PD_H[2]:I PD_H_I2C:I TIE_LO_ESD:O VCC_IO:I
*.PININFO VGND_IO:I
XI97 PD_H[3] net80 sky130_fd_io__tk_em2s
XI108 PD_H[3] net78 sky130_fd_io__tk_em2s
XI109 TIE_LO_ESD net76 sky130_fd_io__tk_em2s
XI102 PD_H[3] net72 sky130_fd_io__tk_em2s
XI104 PD_H[3] net68 sky130_fd_io__tk_em2s
XI96 PD_H[3] net66 sky130_fd_io__tk_em2s
XI113 PD_H[2] net46 sky130_fd_io__tk_em2s
XI99 TIE_LO_ESD net80 sky130_fd_io__tk_em2o
XI98 PD_H[2] net80 sky130_fd_io__tk_em2o
XI106 PD_H[2] net78 sky130_fd_io__tk_em2o
XI107 TIE_LO_ESD net78 sky130_fd_io__tk_em2o
XI110 PD_H[3] net76 sky130_fd_io__tk_em2o
XI111 PD_H[2] net76 sky130_fd_io__tk_em2o
XI100 TIE_LO_ESD net72 sky130_fd_io__tk_em2o
XI101 PD_H[2] net72 sky130_fd_io__tk_em2o
XI103 TIE_LO_ESD net68 sky130_fd_io__tk_em2o
XI105 PD_H[2] net68 sky130_fd_io__tk_em2o
XI95 PD_H[2] net66 sky130_fd_io__tk_em2o
XI94 TIE_LO_ESD net66 sky130_fd_io__tk_em2o
XI88 PD_H[3] net46 sky130_fd_io__tk_em2o
XI87 TIE_LO_ESD net46 sky130_fd_io__tk_em2o
XI49 VGND_IO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xn24<2>_q0 PAD net80 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1>_q0 PAD net80 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0>_q0 PAD net80 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2>_q0 PAD net66 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1>_q0 PAD net66 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0>_q0 PAD net66 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn12_q0 PAD PD_H_I2C VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2>_q0 PAD net68 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1>_q0 PAD net68 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0>_q0 PAD net68 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2>_q0 PAD net78 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1>_q0 PAD net78 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0>_q0 PAD net78 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn13_q0 PAD net46 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn31_q0 PAD net72 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
xI72 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpiov2_pddrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong DRVLO_H_N I2C_MODE_H_N PD_H[4]
+ PD_H[3] PD_H[2] PDEN_H_N SLOW_H TIE_HI_ESD VCC_IO VGND VGND_IO
*.PININFO DRVLO_H_N:I I2C_MODE_H_N:I PD_H[4]:O PD_H[3]:O PD_H[2]:O
*.PININFO PDEN_H_N:I SLOW_H:I TIE_HI_ESD:I VCC_IO:I VGND:I VGND_IO:I
XI160 I2C_MODE_H_N SLOW_H net75 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI98 i2c_mode_h SLOW_H int_slow1 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI161 net75 net142 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI97 int_slow1 mod_slow_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI93 I2C_MODE_H_N i2c_mode_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xmux_q0 mod_drvlo_h_n_i2c DRVLO_H_N i2c_mode_h I2C_MODE_H_N VCC_IO VGND_IO
+ mod_drvlo_h_n sky130_fd_io__gpiov2_octl_mux
Xnr3_q0 DRVLO_H_N pbias_out pbias_out mod_slow_h PD_H[2] PD_H[4] PDEN_H_N VCC_IO
+ VGND_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
Xnr2_q0 mod_drvlo_h_n en_fast2_n<1> en_fast2_n<0> mod_slow_h PD_H[3] PDEN_H_N
+ VCC_IO VGND_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI76 net118 pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> VCC_IO sky130_fd_io__tk_opti
Xinv_q0 en_fast_h en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xbias_q0 DRVLO_H_N en_fast_h en_fast_h_n pbias_out PD_H[4] PDEN_H_N VCC_IO
+ VGND_IO sky130_fd_io__com_pdpredrvr_pbias
Xnor_q0 net142 PDEN_H_N en_fast_h VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI87 mod_drvlo_h_n_i2c PD_H[4] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI88 mod_drvlo_h_n_i2c PD_H[4] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pdpredrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] I2C_MODE_H PD_H PD_I2C_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I I2C_MODE_H:I
*.PININFO PD_H:O PD_I2C_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
Xmpin_slow_q0 PD_I2C_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_I2C_H DRVLO_H_N net62 VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=0.42 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_I2C_H DRVLO_H_N net62 VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=0.42 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast1_q0 net62 EN_FAST_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI72<1> net53<0> EN_FAST_N[1] net42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI72<0> net53<1> EN_FAST_N[0] net42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI74<1> PD_H DRVLO_H_N net53<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74<0> PD_H DRVLO_H_N net53<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI75 net039 PDEN_H_N net42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI76 PD_H DRVLO_H_N net45 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI73 net42 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI101 net45 PDEN_H_N net039 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI94 PD_H I2C_MODE_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnin_q0 PD_I2C_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2
+ w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_q0 PD_I2C_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI78 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pdpredrvr_strong_nr2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] I2C_MODE_H PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I I2C_MODE_H:I
*.PININFO PD_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
XI85 int1 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_slow_q0 PD_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=2.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_H DRVLO_H_N int_nor<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_H DRVLO_H_N int_nor<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast<1>_q0 int_nor<1> EN_FAST_N[1] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_fast<0>_q0 int_nor<0> EN_FAST_N[0] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI90 PD_H DRVLO_H_N net43 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 net43 PDEN_H_N int1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI87<1> PD_H DRVLO_H_N int2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI87<0> PD_H DRVLO_H_N int2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI86<1> int2 EN_FAST_N[1] int1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI86<0> int2 EN_FAST_N[0] int1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnin_q0 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnen_q0 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pdpredrvr_strong_nr3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong DRVHI_H PU_H_N[3] PU_H_N[2] PUEN_H
+ SLOW_H_N VCC_IO VGND_IO
*.PININFO DRVHI_H:I PU_H_N[3]:O PU_H_N[2]:O PUEN_H:I SLOW_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xnd2b_q0 DRVHI_H en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0>
+ PU_H_N[3] PUEN_H VCC_IO VGND_IO sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xnd2a_q0 DRVHI_H net54 net54 net54 net54 PU_H_N[2] PUEN_H VCC_IO VGND_IO
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h sky130_fd_io__tk_opto
Xinv_q0 en_fast_h_n en_fast_h VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xnbias_q0 DRVHI_H en_fast_h en_fast_h_n nbias_out PU_H_N[2] PUEN_H VCC_IO
+ VGND_IO sky130_fd_io__com_pupredrvr_nbias
Xnand_q0 PUEN_H SLOW_H_N en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
.ENDS sky130_fd_io__gpiov2_pupredrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong_nd2 DRVHI_H EN_FAST[3] EN_FAST[2]
+ EN_FAST[1] EN_FAST[0] PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_FAST[3]:I EN_FAST[2]:I EN_FAST[1]:I
*.PININFO EN_FAST[0]:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XE1 net24 PU_H_N sky130_fd_io__tk_em1s
XRrespu1 int_res net24 sky130_fd_pr__res_generic_po W=0.33 L=11 m=1
XRrespu2 PU_H_N int_res sky130_fd_pr__res_generic_po W=0.33 L=4 m=1
Xmnin_fast<3>_q0 net24 DRVHI_H int<3> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<2>_q0 net24 DRVHI_H int<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<1>_q0 net24 DRVHI_H int<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<0>_q0 net24 DRVHI_H int<0> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_slow1_q0 n<2> PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_slow_q0 PU_H_N DRVHI_H n<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_fast<3>_q0 int<3> EN_FAST[3] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<2>_q0 int<2> EN_FAST[2] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<1>_q0 int<1> EN_FAST[1] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<0>_q0 int<0> EN_FAST[0] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_q0 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_q0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pupredrvr_strong_nd2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf IN_H MODE_VCCHIB_LV_N OUT OUT_N
+ VCCHIB VSSD
*.PININFO IN_H:I MODE_VCCHIB_LV_N:I OUT:O OUT_N:O VCCHIB:I VSSD:I
XI420 net57 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI552 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI544 fbk IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI551 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI424 net81 in_b VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI423 OUT_N net81 VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI545 in_b IN_H fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI487 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 m=3 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI541 net81 MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI549 net57 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI436 net81 in_b net112 VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI543 in_b IN_H net108 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI429 OUT_N net81 VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI538 net112 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI489 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI547 net108 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=3 w=5.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_vcchib_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x1 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x2 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x4 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x8 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_nand2 IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_nand2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_nor IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net16 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net16 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_nor

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_xor IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net29 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT net54 net45 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 net70 IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 net54 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 net45 IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT net70 net29 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net58 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net70 IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT net70 net62 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net62 net54 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 net58 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 net54 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_xor

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__inv_1 A Y VGND VNB VPB VPWR
*.PININFO A:I Y:O VGND:I VNB:I VPB:I VPWR:I
XMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__inv_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nand2_1 A B Y VGND VNB VPB VPWR
*.PININFO A:I B:I Y:O VGND:I VNB:I VPB:I VPWR:I
XMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nand2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nand2_2_enhpath IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nand2_2_enhpath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nor2_1 A B Y VGND VNB VPB VPWR
*.PININFO A:I B:I Y:O VGND:I VNB:I VPB:I VPWR:I
XMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nor2_4_enhpath IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net16 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net16 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nor2_4_enhpath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nor3_dnw IN0 IN1 IN2 OUT VGND VPWR
*.PININFO IN0:I IN1:I IN2:I OUT:O VGND:I VPWR:I
XI3 net43 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net39 IN1 net43 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 OUT IN2 net39 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 OUT IN2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nor3_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__res250only_small PAD ROUT
*.PININFO PAD:B ROUT:B

* NOTE: Removed all but the primary resistor;  the other devices do not
* show up in the layout.
*
* RI175 net12 net16 sky130_fd_pr__res_generic_po W=2 L=10.07 m=1
* RI229 net16 ROUT sky130_fd_pr__res_generic_po W=2 L=0.17 m=1
* RI228 PAD net12 sky130_fd_pr__res_generic_po W=2 L=0.17 m=1
* RI237<1> net16 ROUT short
* RI237<2> net16 ROUT short
* RI234<1> PAD net12 short
* RI234<2> PAD net12 short

XRI175 PAD ROUT sky130_fd_pr__res_generic_po W=2 L=10.07 m=1
.ENDS sky130_fd_io__res250only_small

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__res75only_small PAD ROUT
*.PININFO PAD:B ROUT:B
XRI175 PAD ROUT sky130_fd_pr__res_generic_po W=2 L=3.15 m=1
.ENDS sky130_fd_io__res75only_small

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  The resistors here are in an annular shape, and they overlap
* between cells such that the center of the resistor connects between the two
* devices.  To be correct, these two nets must come out as pins.

.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term GATE IN NBODY NWELLRING VGND net16
*.PININFO GATE:I IN:B NBODY:B NWELLRING:B VGND:B
XI1 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=5.4 l=0.6 mult=1
+ sa=0.0 sb=0.0 sd=0.0 topography=normal area=0.048 perim=0.94
* RI9 net18 NBODY short
* RI8 net16 NWELLRING short
RI9 net18 NBODY sky130_fd_pr__res_generic_m1 W=0.02 L=0.005
RI8 net16 NWELLRING sky130_fd_pr__res_generic_m1 W=0.02 L=0.005
.ENDS sky130_fd_io__signal_5_sym_hv_local_5term

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_dly IN OUT OUT_N VCC_IO VGND
*.PININFO IN:I OUT:O OUT_N:O VCC_IO:I VGND:I
XI228 OUT_N a5 sky130_fd_io__tk_em1o
XI229 OUT_N a7 sky130_fd_io__tk_em1o
XI227 a6 OUT sky130_fd_io__tk_em1o
XI214 OUT_N a1 sky130_fd_io__tk_em1o
XI215 a2 OUT sky130_fd_io__tk_em1o
XEdly0 IN OUT sky130_fd_io__tk_em1o
XI217 OUT_N a3 sky130_fd_io__tk_em1s
XEdly2 a4 OUT sky130_fd_io__tk_em1s
XI196 a1 IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI204 a4 a3 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI199 a2 a1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI198 a3 a2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI232 a5 a4 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI231 a6 a5 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI230 a7 a6 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI197 a1 IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI202 a4 a3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI201 a2 a1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI200 a3 a2 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI235 a5 a4 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI234 a6 a5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI233 a7 a6 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_dly

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_hys IN OUT VCC_IO VGND
*.PININFO IN:I OUT:O VCC_IO:I VGND:I
XI650 vcc_io_buf OUT int_n VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI649 int_n IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI648 OUT IN int_n VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI655 vgnd_buf VCC_IO VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI647 vgnd_buf OUT int_p VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI656 vcc_io_buf VGND VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI646 OUT IN int_p VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI645 int_p IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_hys

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_log_i2c_fix DISHS_H DISHS_H_N EN_H ENHS_H
+ ENHS_H_N ENHS_LAT_H_N EXITHS_H FORCEHI_H[1] OD_I_H_N VCC_IO VGND
*.PININFO DISHS_H:O DISHS_H_N:O EN_H:I ENHS_H:O ENHS_H_N:O
*.PININFO ENHS_LAT_H_N:I EXITHS_H:O FORCEHI_H[1]:I OD_I_H_N:I VCC_IO:I
*.PININFO VGND:I
XI664 net39 net46 DISHS_H VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_nand2
XI663 net80 FORCEHI_H[1] net46 VGND VGND VCC_IO VCC_IO
+ sky130_fd_io__sio_hvsbt_nand2
XI662 OD_I_H_N EN_H net39 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_nand2
XI658 OD_I_H_N net80 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI666 ENHS_LAT_H_N net74 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI565 net74 ENHS_H_N VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI667 DISHS_H DISHS_H_N VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI637 ENHS_H_N ENHS_H VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI553 net74 enhs_dly_h_n EXITHS_H VGND VGND VCC_IO VCC_IO
+ sky130_fd_io__sio_hvsbt_nor
XI521 net74 enhs_dly_h enhs_dly_h_n VCC_IO VGND sky130_fd_io__sio_hotswap_dly
.ENDS sky130_fd_io__sio_hotswap_log_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_pghspd IN1 IN2 OUT VGND
*.PININFO IN1:I IN2:I OUT:O VGND:I
XEin2b VGND net25 sky130_fd_io__tk_em1o
XEoutb net38 OUT sky130_fd_io__tk_em1o
XEin1b VGND net27 sky130_fd_io__tk_em1o
XEin1a IN1 net27 sky130_fd_io__tk_em1s
XEouta net42 OUT sky130_fd_io__tk_em1s
XEin2a IN2 net25 sky130_fd_io__tk_em1s
XI481 net50 IN2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI507 OUT IN1 net50 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI651 net42 net27 net34 VGND sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI654 net38 net27 net30 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI652 net34 net25 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI653 net30 net25 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_pghspd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_wpd E_N OUT VGND
*.PININFO E_N:I OUT:O VGND:I
XI198 npd<15> npd<16> sky130_fd_io__tk_em1o
XI209 VGND npd<14> sky130_fd_io__tk_em1o
XI196 npd<17> npd<18> sky130_fd_io__tk_em1o
XI197 npd<16> npd<17> sky130_fd_io__tk_em1o
XE20 npd<18> OUT sky130_fd_io__tk_em1o
XI208 npd<14> npd<15> sky130_fd_io__tk_em1o
Xnen17_q0 npd<17> E_N npd<16> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen15_q0 npd<15> E_N npd<14> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen14_q0 npd<14> E_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen16_q0 npd<16> E_N npd<15> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen19_q0 OUT E_N npd<18> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen18_q0 npd<18> E_N npd<17> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_wpd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x1 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_inv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x2 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_inv_x2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x4 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_inv_x4

.SUBCKT sky130_fd_io__gpio_ovtv2_hvsbt_inv_x4 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_hvsbt_inv_x4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_nand2 IN0 IN1 OUT VGND VNB VPB VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI3 OUT IN0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_nand2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_nor IN0 IN1 OUT VGND VNB VPB VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI3 net17 IN0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net17 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_nor

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_tk_em1o A B
*.PININFO A:B B:B
* RI1 A net11 short
* RI2 B net7 short
RI1 A net11 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI2 B net7 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__sio_tk_em1o

.SUBCKT sky130_fd_io__sio_tk_em2o A B
*.PININFO A:B B:B
RI1 A net11 sky130_fd_pr__res_generic_m2 W=0.66 L=0.01
RI2 B net7 sky130_fd_pr__res_generic_m2 W=0.66 L=0.01
.ENDS sky130_fd_io__sio_tk_em2o

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_tk_em1s A B
*.PININFO A:B B:B
* RI1 A net8 short
* RI2 B net8 short
RI1 A net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI2 B net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__sio_tk_em1s

.SUBCKT sky130_fd_io__sio_tk_em2s A B
*.PININFO A:B B:B
RI1 A net8 sky130_fd_pr__res_generic_m2 W=0.66 L=0.01
RI2 B net8 sky130_fd_pr__res_generic_m2 W=0.66 L=0.01
.ENDS sky130_fd_io__sio_tk_em2s

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_tk_tie_r_out_esd A B
*.PININFO A:B B:B
XResd_r A B sky130_fd_pr__res_generic_po W=0.5 L=10.2 m=1
.ENDS sky130_fd_io__sio_tk_tie_r_out_esd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em1o A B
*.PININFO A:B B:B
* RI1 A net11 short
* RI2 B net7 short
RI1 A net11 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI2 B net7 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__tk_em1o


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em1s A B
*.PININFO A:B B:B
* RI1 A net8 short
* RI2 B net8 short
RI1 A net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI2 B net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__tk_em1s


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em2o A B
*.PININFO A:B B:B
* RI1 A net11 short
* RI2 B net7 short
RI1 A net11 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
RI2 B net7 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
.ENDS sky130_fd_io__tk_em2o

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em2s A B
*.PININFO A:B B:B
* RI1 A net8 short
* RI2 B net8 short
RI1 A net8 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
RI2 B net8 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
.ENDS sky130_fd_io__tk_em2s

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_opti OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em1o
Xe1_q0 OUT SPU sky130_fd_io__tk_em1s
.ENDS sky130_fd_io__tk_opti


* optiA is the same as opti, but uses tk_em2s, which is like tk_em1s
* but with a m2 short instead of a m1 short.

.SUBCKT sky130_fd_io__tk_optiA OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em1o
Xe1_q0 OUT SPU sky130_fd_io__tk_em2s
.ENDS sky130_fd_io__tk_optiA

* optiB is the same as opti, but uses tk_em2s, which is like tk_em1s
* but with a m2 short instead of a m1 short, and tk_em2o, which is
* like tk_em1o but with m2 shorts instead of m1 shorts.

.SUBCKT sky130_fd_io__tk_optiB OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em2o
Xe1_q0 OUT SPU sky130_fd_io__tk_em2s
.ENDS sky130_fd_io__tk_optiB

* optiC is the same as opti, but uses tk_em2o, which is like tk_em1o
* but with an m2 open instead of an m1 open.

.SUBCKT sky130_fd_io__tk_optiC OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em2o
Xe1_q0 OUT SPU sky130_fd_io__tk_em1s
.ENDS sky130_fd_io__tk_optiC

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_opto OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe1_q0 SPU OUT sky130_fd_io__tk_em1o
Xe2_q0 OUT SPD sky130_fd_io__tk_em1s
.ENDS sky130_fd_io__tk_opto

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_tie_r_out_esd A B
*.PININFO A:B B:B
XResd_r A B sky130_fd_pr__res_generic_po W=0.5 L=10.2 m=1
.ENDS sky130_fd_io__tk_tie_r_out_esd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_amuxsplitv2 AMUXBUS_A_L AMUXBUS_A_R AMUXBUS_B_L
+ AMUXBUS_B_R ENABLE_VDDA_H HLD_VDDA_H_N SWITCH_AA_S0 SWITCH_AA_SL SWITCH_AA_SR
+ SWITCH_BB_S0 SWITCH_BB_SL SWITCH_BB_SR VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD
+ VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A_L:B AMUXBUS_A_R:B AMUXBUS_B_L:B AMUXBUS_B_R:B
*.PININFO ENABLE_VDDA_H:I HLD_VDDA_H_N:I SWITCH_AA_S0:I SWITCH_AA_SL:I
*.PININFO SWITCH_AA_SR:I SWITCH_BB_S0:I SWITCH_BB_SL:I SWITCH_BB_SR:I
*.PININFO VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B VSSA:B VSSD:B
*.PININFO VSSIO:B VSSIO_Q:B VSWITCH:B
xI22 VSSA VDDA sky130_fd_io__condiode
XI18 hold SWITCH_AA_S0 ng_vdda_aa_s0_h reset VCCD VDDA VSSA VSSD
+ sky130_fd_io__amuxsplitv2_switch_s0
XI348 hold SWITCH_BB_S0 ng_vdda_bb_s0_h reset VCCD VDDA VSSA VSSD
+ sky130_fd_io__amuxsplitv2_switch_s0
XI347 hold SWITCH_AA_SL ng_vswitch_aa_sl_h pg_vdda_aa_sl_h_n reset VCCD VDDA
+ VSSA VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI24 hold SWITCH_AA_SR ng_vswitch_aa_sr_h pg_vdda_aa_sr_h_n reset VCCD VDDA VSSA
+ VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI349 hold SWITCH_BB_SR ng_vswitch_bb_sr_h pg_vdda_bb_sr_h_n reset VCCD VDDA
+ VSSA VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI350 hold SWITCH_BB_SL ng_vswitch_bb_sl_h pg_vdda_bb_sl_h_n reset VCCD VDDA
+ VSSA VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI6 AMUXBUS_A_L AMUXBUS_A_R ng_vswitch_aa_sl_h ng_vswitch_aa_sr_h
+ ng_vdda_aa_s0_h pg_vdda_aa_sl_h_n pg_vdda_aa_sr_h_n VDDA VSSA
+ sky130_fd_io__amuxsplitv2_switch
XI8 AMUXBUS_B_L AMUXBUS_B_R ng_vswitch_bb_sl_h ng_vswitch_bb_sr_h
+ ng_vdda_bb_s0_h pg_vdda_bb_sl_h_n pg_vdda_bb_sr_h_n VDDA VSSA
+ sky130_fd_io__amuxsplitv2_switch
XI342 ENABLE_VDDA_H HLD_VDDA_H_N hold reset VDDA VSSA
+ sky130_fd_io__amuxsplitv2_delay
.ENDS sky130_fd_io__top_amuxsplitv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_gpio_ovtv2 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL
+ ANALOG_SEL DM[2] DM[1] DM[0] ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO
+ ENABLE_VSWITCH_H HLD_H_N HLD_OVR HYS_TRIM IB_MODE_SEL[1] IB_MODE_SEL[0] IN IN_H
+ INP_DIS OE_N OUT PAD PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H SLEW_CTL[1]
+ SLEW_CTL[0] SLOW TIE_HI_ESD TIE_LO_ESD VCCD VCCHIB VDDA VDDIO VDDIO_Q VINREF
+ VSSA VSSD VSSIO VSSIO_Q VSWITCH VTRIP_SEL
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I DM[2]:I DM[1]:I DM[0]:I ENABLE_H:I
*.PININFO ENABLE_INP_H:I ENABLE_VDDA_H:I ENABLE_VDDIO:I
*.PININFO ENABLE_VSWITCH_H:I HLD_H_N:I HLD_OVR:I HYS_TRIM:I
*.PININFO IB_MODE_SEL[1]:I IB_MODE_SEL[0]:I IN:O IN_H:O INP_DIS:I
*.PININFO OE_N:I OUT:I PAD:B PAD_A_ESD_0_H:B PAD_A_ESD_1_H:B
*.PININFO PAD_A_NOESD_H:B SLEW_CTL[1]:I SLEW_CTL[0]:I SLOW:I
*.PININFO TIE_HI_ESD:O TIE_LO_ESD:O VCCD:B VCCHIB:B VDDA:B VDDIO:B
*.PININFO VDDIO_Q:B VINREF:I VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
*.PININFO VTRIP_SEL:I
Xopath_q0 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n
+ hld_i_ovr_h nga_pad_vpmp_h ngb_pad_vpmp_h od_i_h_n OE_N OUT PAD pd_csd_h pghs_h
+ pu_csd_h pug_h<6> pug_h<5> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1>
+ slew_ctl_h_n<0> SLOW TIE_HI_ESD TIE_LO_ESD VCCD VDDIO VDDIO_Q vpb_drvr VCCHIB
+ VSSA VSSD VSSIO VSSIO_Q sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix
Xovt_amux_q0 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H
+ ENABLE_VSWITCH_H hld_i_h_n nga_pad_vpmp_h ngb_pad_vpmp_h TIE_HI_ESD OUT PAD
+ pd_csd_h pghs_h pu_csd_h pug_h<6> pug_h<5> VCCD VDDA VDDIO VDDIO_Q vpb_drvr VSSA
+ VSSD VSSIO VSWITCH sky130_fd_io__gpio_ovtv2_amux_i2c_fix
Xctrl_q0 DM[2] DM[1] DM[0] dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0>
+ ENABLE_H ENABLE_INP_H HLD_H_N hld_i_h_n hld_i_ovr_h HLD_OVR HYS_TRIM hyst_trim_h
+ net164 IB_MODE_SEL[1] IB_MODE_SEL[0] ib_mode_sel_h<1> ib_mode_sel_h<0> net166<0>
+ net166<1> INP_DIS inp_dis_h_n od_i_h_n SLEW_CTL[1] SLEW_CTL[0] slew_ctl_h<1>
+ slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> VCCD VDDIO_Q VSSD VTRIP_SEL
+ vtrip_sel_h sky130_fd_io__gpio_ctlv2_i2c_fix
XI336 net193 PAD_A_ESD_1_H sky130_fd_io__res75only_small
XI335 PAD net193 sky130_fd_io__res75only_small
XI334 net189 PAD_A_ESD_0_H sky130_fd_io__res75only_small
Xresd4_q0 PAD net189 sky130_fd_io__res75only_small
Xipath_q0 dm_h_n<2> dm_h_n<1> dm_h_n<0> ENABLE_VDDIO hyst_trim_h
+ ib_mode_sel_h<1> ib_mode_sel_h<0> inp_dis_h_n IN IN_H PAD VCCHIB VDDIO_Q VINREF
+ VSSD vtrip_sel_h sky130_fd_io__gpio_ovtv2_ipath
* RS0 PAD PAD_A_NOESD_H short
RS0 PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m4 W=0.88 L=0.01
.ENDS sky130_fd_io__top_gpio_ovtv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_gpiov2 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL
+ ANALOG_SEL DM[2] DM[1] DM[0] ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO
+ ENABLE_VSWITCH_H HLD_H_N HLD_OVR IB_MODE_SEL IN IN_H INP_DIS OE_N OUT PAD
+ PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H SLOW TIE_HI_ESD TIE_LO_ESD VCCD VCCHIB
+ VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH VTRIP_SEL
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I DM[2]:I DM[1]:I DM[0]:I ENABLE_H:I
*.PININFO ENABLE_INP_H:I ENABLE_VDDA_H:I ENABLE_VDDIO:I
*.PININFO ENABLE_VSWITCH_H:I HLD_H_N:I HLD_OVR:I IB_MODE_SEL:I IN:O
*.PININFO IN_H:O INP_DIS:I OE_N:I OUT:I PAD:B PAD_A_ESD_0_H:B
*.PININFO PAD_A_ESD_1_H:B PAD_A_NOESD_H:B SLOW:I TIE_HI_ESD:O
*.PININFO TIE_LO_ESD:O VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B VSSA:B
*.PININFO VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B VTRIP_SEL:I
Xamux_q0 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H
+ ENABLE_VSWITCH_H hld_i_h hld_i_h_n OUT PAD VCCD VDDA VDDIO_Q VSSA VSSD VSSIO_Q
+ VSWITCH sky130_fd_io__gpiov2_amux
Xopath_q0 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n
+ hld_i_ovr_h od_i_h OE_N OUT PAD SLOW TIE_HI_ESD TIE_LO_ESD VDDIO VSSD VSSIO VCCD
+ VCCHIB sky130_fd_io__gpiov2_opath
Xctrl_q0 DM[2] DM[1] DM[0] dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0>
+ ENABLE_H ENABLE_INP_H HLD_H_N hld_i_h hld_i_h_n hld_i_ovr_h HLD_OVR IB_MODE_SEL
+ ib_mode_sel_h ib_mode_sel_h_n INP_DIS inp_dis_h_n od_i_h VDDIO_Q VSSD VCCD
+ VTRIP_SEL vtrip_sel_h vtrip_sel_h_n sky130_fd_io__gpiov2_ctl
Xipath_q0 dm_h_n<2> dm_h_n<1> dm_h_n<0> ENABLE_VDDIO ib_mode_sel_h
+ ib_mode_sel_h_n inp_dis_h_n IN IN_H PAD VCCHIB VDDIO_Q VSSD vtrip_sel_h_n
+ sky130_fd_io__gpiov2_ipath
Xresd3_q0 PAD_A_ESD_1_H net210 sky130_fd_io__res75only_small
Xresd1_q0 net204 PAD sky130_fd_io__res75only_small
Xresd4_q0 net210 PAD sky130_fd_io__res75only_small
Xresd2_q0 PAD_A_ESD_0_H net204 sky130_fd_io__res75only_small
* RS0<2> PAD PAD_A_NOESD_H short
* RS0<1> PAD PAD_A_NOESD_H short
* RS0<0> PAD PAD_A_NOESD_H short
RS0<2> PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m4 W=12.35 L=0.035
RS0<1> PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m3 W=1.07 L=0.035
RS0<0> PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m3 W=12.37 L=0.035
.ENDS sky130_fd_io__top_gpiov2


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_ground_hvc_wpad AMUXBUS_A AMUXBUS_B DRN_HVC G_CORE
+ G_PAD OGC_HVC PADISOL PADISOR SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA
+ VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B DRN_HVC:B G_CORE:B G_PAD:B OGC_HVC:B
*.PININFO PADISOL:B PADISOR:B SRC_BDY_HVC:B VCCD:B VCCHIB:B VDDA:B VDDIO:B
*.PININFO VDDIO_L:B VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
xI39 SRC_BDY_HVC VDDIO sky130_fd_io__condiode
Xcxtor2_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=22 w=10.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc2_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=5 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc1_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xpre_n1_q0 g_nclamp g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xclamp_xtor_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC
+ sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XRrc_res g_pdpre net94 sky130_fd_pr__res_generic_po W=0.33 L=470 m=1
XRI38 net90 DRN_HVC sky130_fd_pr__res_generic_po W=0.33 L=700 m=1
XRI37 net94 net90 sky130_fd_pr__res_generic_po W=0.33 L=1550 m=1
Xpre_p1_q0 g_nclamp g_pdpre DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 m=50
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
RI13 G_PAD G_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
.ENDS sky130_fd_io__top_ground_hvc_wpad

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_hvclampv2 DRN_HVC OGC_HVC SRC_BDY_HVC VSSD
*.PININFO DRN_HVC:B OGC_HVC:B SRC_BDY_HVC:B VSSD:B
xI39 SRC_BDY_HVC OGC_HVC sky130_fd_io__condiode
Xpre_p1_q0 g_nclamp g_pdpre DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 m=50
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XRrc_res g_pdpre net41 sky130_fd_pr__res_generic_po W=0.33 L=470 m=1
XRI38 net37 DRN_HVC sky130_fd_pr__res_generic_po W=0.33 L=700 m=1
XRI37 net41 net37 sky130_fd_pr__res_generic_po W=0.33 L=1550 m=1
Xclamp_xtor_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC
+ sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc1_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc2_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=5 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xcxtor2_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=22 w=10.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__top_hvclampv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 AMUXBUS_A AMUXBUS_B DRN_HVC OGC_HVC
+ PADISOL PADISOR P_CORE P_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA
+ VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B DRN_HVC:B OGC_HVC:B PADISOL:B PADISOR:B
*.PININFO P_CORE:B P_PAD:B SRC_BDY_HVC:B VCCD:B VCCHIB:B VDDA:B VDDIO:B
*.PINFNFO VDDIO_Q:B VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
xI39 SRC_BDY_HVC VDDIO sky130_fd_io__condiode
Xpre_p1_q0 g_nclamp g_pdpre DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 m=50
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XRrc_res g_pdpre net67 sky130_fd_pr__res_generic_po W=0.33 L=470 m=1
XRI38 net63 DRN_HVC sky130_fd_pr__res_generic_po W=0.33 L=700 m=1
XRI37 net67 net63 sky130_fd_pr__res_generic_po W=0.33 L=1550 m=1
Xclamp_xtor_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC
+ sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc1_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc2_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=5 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xcxtor2_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=22 w=10.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
RI13 P_PAD P_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL P_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR P_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
.ENDS sky130_fd_io__top_power_hvc_wpadv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_vrefcapv2 AMUXBUS_A AMUXBUS_B CNEG CPOS VCCD VCCHIB
+ VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B CNEG:B CPOS:B VCCD:B VCCHIB:B VDDA:B
*.PININFO VDDIO:B VDDIO_Q:B VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
xI271 CNEG VDDIO_Q sky130_fd_io__condiode
XI334 CNEG CPOS CNEG CNEG sky130_fd_pr__nfet_05v0_nvt m=180 w=10.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__top_vrefcapv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  Split power and ground nets on XI364<1:0> fixed

.SUBCKT sky130_fd_io__top_xres4v2 AMUXBUS_A AMUXBUS_B DISABLE_PULLUP_H
+ EN_VDDIO_SIG_H ENABLE_H ENABLE_VDDIO FILT_IN_H INP_SEL_H PAD PAD_A_ESD_H
+ PULLUP_H TIE_HI_ESD TIE_LO_ESD TIE_WEAK_HI_H VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA
+ VSSD VSSIO VSSIO_Q VSWITCH XRES_H_N
*.PININFO AMUXBUS_A:B AMUXBUS_B:B DISABLE_PULLUP_H:I EN_VDDIO_SIG_H:I
*.PININFO ENABLE_H:I ENABLE_VDDIO:I FILT_IN_H:I INP_SEL_H:I PAD:B
*.PININFO PAD_A_ESD_H:B PULLUP_H:B TIE_HI_ESD:O TIE_LO_ESD:O
*.PININFO TIE_WEAK_HI_H:B VCCD:I VCCHIB:I VDDA:I VDDIO:I VDDIO_Q:I
*.PININFO VSSA:I VSSD:I VSSIO:I VSSIO_Q:I VSWITCH:I XRES_H_N:O
XI326 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
XI49 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xgpio_inbuf_q0 ENABLE_H ENABLE_VDDIO net79 net83 in_h VCCHIB VDDIO_Q VSSD
+ EN_VDDIO_SIG_H en_vddio_sig_h_n sky130_fd_io__xres4v2_in_buf
Xxresesd_q0 in_h net86 PAD VDDIO VSSD VSSIO sky130_fd_io__xres_esd
Xweakpullup_q0 TIE_WEAK_HI_H VDDIO VSSD sky130_fd_io__xres_wpu
Xesd_res_q0 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
XI335 net97 PULLUP_H VSSD sky130_fd_io__com_xres_weak_pu
XI363 INP_SEL_H inp_sel_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x2
XI334 net103 net107 VSSD VDDIO sky130_fd_io__hvsbt_inv_x2
XI333 DISABLE_PULLUP_H net103 VSSD VDDIO sky130_fd_io__hvsbt_inv_x2
XI374 EN_VDDIO_SIG_H en_vddio_sig_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x2
XI368 net124 out_rcfilt_h VDDIO_Q VSSD sky130_fd_io__xres_rcfilter_lpf
XI367 out_rcfilt_h out_hysbuf_h VDDIO_Q VSSD sky130_fd_io__xres_inv_hys
XI365 out_hysbuf_h out_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI364<1> out_h_n XRES_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x4
XI364<0> out_h_n XRES_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x4
XI361 net124 inp_sel_h_n FILT_IN_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI358 net124 INP_SEL_H net79 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI332 net97 net107 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI360 net124 INP_SEL_H FILT_IN_H VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI357 net124 inp_sel_h_n net79 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__top_xres4v2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xor2_1 A B X VGND VPWR
*.PININFO A:I B:I X:O VGND:I VPWR:I
XMNnor0 inor A VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNnor1 inor B VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNaoi10 VGND A sndNA VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNaoi11 sndNA B X VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNaoi20 X inor VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPnor0 VPWR A sndPA VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPnor1 sndPA B inor VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPaoi10 pmid A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPaoi11 pmid B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPaoi20 X inor pmid VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres4v2_in_buf ENABLE_HV ENABLE_VDDIO_LV IN_H IN_H_N PAD
+ VCCHIB VDDIO VGND VNORMAL VNORMAL_B
*.PININFO ENABLE_HV:I ENABLE_VDDIO_LV:I IN_H:O IN_H_N:O PAD:I VCCHIB:I
*.PININFO VDDIO:I VGND:I VNORMAL:I VNORMAL_B:I
XI165 ENABLE_VDDIO_LV enable_vddio_lv_n VGND VGND VCCHIB VCCHIB
+ sky130_fd_io__inv_1
XI61 net106 mode_vcchib VGND VDDIO sky130_fd_io__hvsbt_inv_x1
XI35 VNORMAL_B ENABLE_HV net106 VGND VDDIO sky130_fd_io__hvsbt_nand2
XI132 net207 net110 VGND sky130_fd_pr__res_generic_nd__hv W=0.29 L=1077.19 m=1
XRI159 net235 net108 sky130_fd_pr__res_generic_po W=0.4 L=713.695 m=1
XI8 net193 pad1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI86 pad1 pad_inv VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85 pad_inv PAD net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI114 net152 pad_inv net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI145 enable_hv_b ENABLE_HV VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI251 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI83 net140 PAD VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 fbk pad_inv VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI213 IN_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI152 VGND VGND VGND VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI113 net124 PAD net152 VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI154 net120 mode_vcchib net206 VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI151 net116 mode_vcchib vcchib_int VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0
+ l=0.9 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI150 net112 pad_inv net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI116 pad1 pad_inv net235 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI143 net124 VNORMAL VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI156 net116 enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI252 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI107 net108 mode_vcchib VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI146 enable_hv_b ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI88 pad_inv PAD vcchib_int vcchib_int sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0
+ l=0.8 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI89 pad_inv PAD net207 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI90 pad1 pad_inv net206 net206 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI133 net110 mode_vcchib VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 net193 fbk VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI219 fbk net193 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 IN_H_N fbk VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI158 net120 enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI139 net207 VNORMAL_B net110 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI136 net112 VNORMAL_B VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI153 vcchib_int vcchib_int vcchib_int vcchib_int sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=1.0 l=0.8 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI160 net235 VNORMAL_B net108 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xres4v2_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_esd OUT_H OUT_VT PAD VDDIO VSSD VSSIO
*.PININFO OUT_H:B OUT_VT:B PAD:B VDDIO:B VSSD:B VSSIO:B
Xesd_q0 PAD OUT_H OUT_VT VDDIO VSSD VSSD sky130_fd_io__gpio_buf_localesd
Xpddrvr_strong_q0 tie_lo_esd tie_lo_esd PAD tie_lo_esd tie_lo_esd tie_lo_esd
+ VDDIO VSSIO VSSIO sky130_fd_io__gpio_pddrvr_strong
Xpudrvr_strong_q0 PAD tie_hi_esd tie_hi_esd tie_hi_esd VDDIO VSSD
+ sky130_fd_io__gpio_pudrvr_strong
xI271 VSSIO VDDIO sky130_fd_io__condiode
.ENDS sky130_fd_io__xres_esd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_inv_hys IN_H OUT_H VCC_IO VSSD
*.PININFO IN_H:I OUT_H:O VCC_IO:I VSSD:I
XI7 pmid1 IN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 out_h_n IN_H pmid1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H out_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI10 pmid1 OUT_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 out_h_n IN_H nmid1 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 nmid1 IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT_H out_h_n VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 nmid1 OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xres_inv_hys

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_rcfilter_lpf IN OUT VCC_IO VSSD
*.PININFO IN:I OUT:O VCC_IO:B VSSD:B
Xe5_q0 net65 net40 sky130_fd_io__xres_tk_emlo
Xe1_q0 net135 net67 sky130_fd_io__xres_tk_emlo
Xe4_q0 net43 net65 sky130_fd_io__xres_tk_emlo
XI200 net59 OUT sky130_fd_io__xres_tk_emlo
XI199 net62 OUT sky130_fd_io__xres_tk_emlo
XI198 VSSD net59 sky130_fd_io__xres_tk_emlo
XI197 VSSD net57 sky130_fd_io__xres_tk_emlo
XI194 net57 OUT sky130_fd_io__xres_tk_emlo
XI193 net45 OUT sky130_fd_io__xres_tk_emlo
XI191 net42 OUT sky130_fd_io__xres_tk_emlo
XI190 net40 OUT sky130_fd_io__xres_tk_emlo
XI187 VSSD OUT sky130_fd_io__xres_tk_emlo
XI186 VSSD net45 sky130_fd_io__xres_tk_emlo
Xe2_q0 net67 net43 sky130_fd_io__xres_tk_emlo
XI183 net42 VSSD sky130_fd_io__xres_tk_emlo
XI181 net40 VSSD sky130_fd_io__xres_tk_emlo
XI202 VSSD sky130_fd_io__xres_tk_emlc
XI201 VSSD sky130_fd_io__xres_tk_emlc
XI192 OUT sky130_fd_io__xres_tk_emlc
XI189 VSSD sky130_fd_io__xres_tk_emlc
XI188 VSSD sky130_fd_io__xres_tk_emlc
XI180 net40 sky130_fd_io__xres_tk_emlc
XI182 net42 sky130_fd_io__xres_tk_emlc
Xe3_q0 net43 sky130_fd_io__xres_tk_emlc
XI172 IN net135 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI184 VSSD net57 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI185 VSSD net45 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI196 VSSD net62 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI195 VSSD net59 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI179 net43 net65 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI178 net65 net40 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI177 net40 net42 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI176 net42 OUT VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI175 net67 net43 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI174 net43 net43 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI173 net135 net67 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
.ENDS sky130_fd_io__xres_rcfilter_lpf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_rcfilter_lpf_rcunit IN OUT VGND VNB VPWR
*.PININFO IN:I OUT:O VGND:B VNB:B VPWR:B
Xr1b_q0 net14 OUT VNB sky130_fd_io__xres_rcfilter_lpf_res_sub
Xr1a_q0 IN net14 VNB sky130_fd_io__xres_rcfilter_lpf_res_sub
XI242 VGND OUT VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=7.0 l=4.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI244 VPWR OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.0 l=4.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xres_rcfilter_lpf_rcunit

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  Added 3rd terminal to sky130_fd_pr__res_generic_nd devices

.SUBCKT sky130_fd_io__xres_rcfilter_lpf_res_sub IN OUT VGND
*.PININFO IN:I OUT:O VGND:B
Xe1_q0 IN sky130_fd_io__xres_tk_emlc
Xe2_q0 OUT net30 sky130_fd_io__xres_tk_emlo
Xropti OUT net30 VGND sky130_fd_pr__res_generic_nd W=0.5 L=14 m=1
Xr1 net30 IN VGND sky130_fd_pr__res_generic_nd W=0.5 L=47 m=1
Xropto IN IN VGND sky130_fd_pr__res_generic_nd W=0.5 L=14 m=1
.ENDS sky130_fd_io__xres_rcfilter_lpf_res_sub

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_tk_emlc A
*.PININFO A:B
* RI2 A net7 short
* RI1 A net2 short
RI2 A net7 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI1 A net2 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__xres_tk_emlc

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_tk_emlo A B
*.PININFO A:B B:B
* RI2 B net8 short
* RI1 A net3 short
RI2 B net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI1 A net3 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__xres_tk_emlo

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_wpu PAD VDDIO VSSD
*.PININFO PAD:B VDDIO:B VSSD:B
Xesdr_q0 PAD net15 sky130_fd_io__res250only_small
X5kres_q0 VDDIO net15 VSSD sky130_fd_io__com_res_weak
.ENDS sky130_fd_io__xres_wpu

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_ground_lvc_wpad AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1
+ DRN_LVC2 G_CORE G_PAD OGC_LVC PADISOL PADISOR SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD
+ VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B BDY2_B2B:B DRN_LVC1:B DRN_LVC2:B
*.PININFO G_CORE:B G_PAD:B OGC_LVC:B PADISOL:B PADISOR:B SRC_BDY_LVC1:B
*.PININFO SRC_BDY_LVC2:B VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B VSSA:B
*.PININFO VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
Xesd_q0 BDY2_B2B SRC_BDY_LVC1 VSSD sky130_fd_io__gnd2gnd_120x2_lv_isosub
xI54 SRC_BDY_LVC2 VDDIO sky130_fd_io__condiode
xI50 SRC_BDY_LVC1 VDDIO sky130_fd_io__condiode
RI21 G_PAD G_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
Xpre_p1_q0 g_nclamp_lvc1 g_pdpre_lvc1 DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8
+ m=20 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI40 g_nclamp_lvc2 g_pdpre_lvc2 DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 m=20
+ w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xclamp_xtor_q0 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=166 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI42 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=152 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI61 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=38 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI62 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8
+ m=20 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xncap_q0 SRC_BDY_LVC1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=15 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp_lvc1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=3 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI43 g_nclamp_lvc2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2
+ sky130_fd_pr__nfet_01v8 m=2 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI58 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=6 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI60 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=1 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI59 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=10 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XRrc_res g_pdpre_lvc1 DRN_LVC1 sky130_fd_pr__res_generic_po W=0.33 L=1950 m=1
XRI44 DRN_LVC2 net161 sky130_fd_pr__res_generic_po W=0.33 L=900 m=1
XRI47 net161 net155 sky130_fd_pr__res_generic_po W=0.33 L=300 m=1
XRI46 g_pdpre_lvc2 net157 sky130_fd_pr__res_generic_po W=0.33 L=200 m=1
XRI45 net157 net155 sky130_fd_pr__res_generic_po W=0.33 L=720 m=1
.ENDS sky130_fd_io__top_ground_lvc_wpad

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_power_lvc_wpad AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1
+ DRN_LVC2 OGC_LVC PADISOL PADISOR P_CORE P_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD
+ VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B BDY2_B2B:B DRN_LVC1:B DRN_LVC2:B
*.PININFO OGC_LVC:B PADISOL:B PADISOR:B P_CORE:B P_PAD:B SRC_BDY_LVC1:B
*.PININFO SRC_BDY_LVC2:B VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B
*.PININFO VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
Xesd_q0 BDY2_B2B SRC_BDY_LVC1 VSSD sky130_fd_io__gnd2gnd_120x2_lv_isosub
xI54 SRC_BDY_LVC2 VDDIO sky130_fd_io__condiode
xI50 SRC_BDY_LVC1 VDDIO sky130_fd_io__condiode
RI21 P_PAD P_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL P_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR P_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
Xpre_p1_q0 g_nclamp_lvc1 g_pdpre_lvc1 DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8
+ m=20 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI40 g_nclamp_lvc2 g_pdpre_lvc2 DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 m=20
+ w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xclamp_xtor_q0 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=166 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI42 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=152 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI61 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=38 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI62 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8
+ m=20 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xncap_q0 SRC_BDY_LVC1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=15 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp_lvc1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=3 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI43 g_nclamp_lvc2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2
+ sky130_fd_pr__nfet_01v8 m=2 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI58 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=6 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI60 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=1 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI59 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=10 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XRrc_res g_pdpre_lvc1 DRN_LVC1 sky130_fd_pr__res_generic_po W=0.33 L=1950 m=1
XRI44 DRN_LVC2 net161 sky130_fd_pr__res_generic_po W=0.33 L=900 m=1
XRI47 net161 net155 sky130_fd_pr__res_generic_po W=0.33 L=300 m=1
XRI46 g_pdpre_lvc2 net157 sky130_fd_pr__res_generic_po W=0.33 L=200 m=1
XRI45 net157 net155 sky130_fd_pr__res_generic_po W=0.33 L=720 m=1
.ENDS sky130_fd_io__top_power_lvc_wpad

* The following subcircuits were added 10/19/2023 and include cells that were
* in earlier versions of the I/O library and which did not get into the first
* build of the sky130_fd_io library.

.SUBCKT sky130_fd_io__top_analog_pad amuxbus_a amuxbus_b pad pad_core vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B pad:B pad_core:B vccd:B vcchib:B vdda:B 
*.PININFO vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
RI289 pad_core pad sky130_fd_pr__res_generic_m3  L=0.9  W=8.98
Xpudrvr_strong pad tie_hi_esd tie_hi_esd tie_hi_esd vddio vssd 
+ sky130_fd_io__gpio_pudrvr_strong
Xpddrvr_strong tie_lo_esd tie_lo_esd pad tie_lo_esd tie_lo_esd tie_lo_esd 
+ vddio vssio vssio sky130_fd_io__gpio_pddrvr_strong
.ENDS

.SUBCKT sky130_fd_io__xres_hvlv_ls in_h out_c out_t vcchib vddio_q vssd
*.PININFO in_h:I vcchib:I vddio_q:I vssd:I out_c:O out_t:O
XI11 in_int_h_n in_int_h vssd vddio_q sky130_fd_io__hvsbt_inv_x1
XI10 in_h in_int_h_n vssd vddio_q sky130_fd_io__hvsbt_inv_x1
XI534 out_t out_c vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_c out_t vcchib vcchib sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI536 out_c in_int_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_t in_int_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__xres_buf_hys in_h out_h vcc_io vssd
*.PININFO in_h:I vcc_io:I vssd:I out_h:O
XI7 pmid1 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 out_h_n in_h pmid1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 out_h out_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 pmid1 out_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 out_h_n in_h nmid1 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 nmid1 in_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 out_h out_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 nmid1 out_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__top_axresv2 amuxbus_a amuxbus_b disable_pullup_h filter_in_h 
+ filter_out filter_out_h pullup_h tie_hi_esd tie_lo_esd vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO disable_pullup_h:I filter_in_h:I filter_out:O filter_out_h:O 
*.PININFO tie_hi_esd:O tie_lo_esd:O amuxbus_a:B amuxbus_b:B pullup_h:B vccd:B 
*.PININFO vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B 
*.PININFO vswitch:B
Xrcfilt filter_in_h out_rcfilt_h vddio_q vssd sky130_fd_io__xres_rcfilter_lpf
Xhv_lv_ls out_hysbuf_h net66 net65 vcchib vddio_q vssd sky130_fd_io__xres_hvlv_ls
Xhv_drv1 out_hysbuf_h out_h_n vssd vddio_q sky130_fd_io__hvsbt_inv_x1
Xhv_drv2 out_h_n filter_out_h vssd vddio_q sky130_fd_io__hvsbt_inv_x4
XI330 net77 pullup_h vssd sky130_fd_io__com_xres_weak_pu
XI323 net86 net93 vssd vddio sky130_fd_io__hvsbt_inv_x2
XI324 disable_pullup_h net86 vssd vddio sky130_fd_io__hvsbt_inv_x2
Xhyst_buf out_rcfilt_h out_hysbuf_h vddio_q vssd sky130_fd_io__xres_buf_hys
XI32 net108 net65 vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI321 net77 net93 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI33 filter_out net108 vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=4 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI326 vssio tie_lo_esd sky130_fd_io__tk_tie_r_out_esd
XI49 vddio tie_hi_esd sky130_fd_io__tk_tie_r_out_esd
XI34 net108 net65 vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI35 filter_out net108 vssd vssd sky130_fd_pr__nfet_01v8 m=8 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_inbuf_lvinv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_inbuf_hvinv_x1 in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_inbuf_hvinv_x2 in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_inbuf_lvinv_x2 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=5.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_in_buf en_h in_h in_vt out_h out_h_n vcc_io vgnd vpwr 
+ vtrip_sel_h_n
*.PININFO en_h:I in_h:I in_vt:I vcc_io:I vgnd:I vpwr:I vtrip_sel_h_n:I out_h:O 
*.PININFO out_h_n:O
XI596 out_a net115 sky130_fd_io__tk_em1s
Xttl_pd_op net077 net118 sky130_fd_io__tk_em1o
XI576 vtrip_sel_h_n vtrip_sel_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xpd2 net134 out_a vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1_mid_nat net130 vpwr net103 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpd_hrng net118 in_vt net117 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=3.00 l=1.00 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpden_1 net117 en_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpd1 net118 in_h net117 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI585 net115 net115 out_a vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI574 net118 out_a net137 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI598 net118 out_a vcc_io vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI592 out_h out_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI584 net103 net103 net115 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI571 net118 out_a vcc_io vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI597 net118 out_a net137 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI570 out_a in_h net118 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI595 net077 in_vt net117 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=3.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI589 out_h_n net134 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xdis_trip_sel1 in_vt vtrip_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu2 net134 out_a vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1 net169 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpuen_2 out_a en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1_midopt net169 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI567 net130 in_h net169 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI568 vgnd out_a net169 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI590 out_h_n net134 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI579 net153 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI578 out_a in_h net153 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI593 out_h out_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI577 out_a vtrip_sel_h net130 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI582 vgnd out_a net153 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI575 vcc_io vtrip_sel_h net137 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__com_ictl_logic analog_en_h dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ inp_dis_h_n inp_dis_i_h inp_dis_i_h_n startup_en_h tripsel_i_h tripsel_i_h_n 
+ vcc_io vgnd vtrip_sel_h
*.PININFO analog_en_h:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I inp_dis_h_n:I 
*.PININFO startup_en_h:I vcc_io:I vgnd:I vtrip_sel_h:I inp_dis_i_h:O 
*.PININFO inp_dis_i_h_n:O tripsel_i_h:O tripsel_i_h_n:O
XI29 net58 analog_en_h net042 vgnd vcc_io sky130_fd_io__hvsbt_nor
XI30 startup_en_h net042 inp_dis_i_h vgnd vcc_io sky130_fd_io__hvsbt_nor
Xinpdis_inv inp_dis_i_h inp_dis_i_h_n vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xdm10nand_inv nand_dm01 and_dm01 vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xtripsel_inv tripsel_i_h_n tripsel_i_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xinpdis dm_buf_dis inp_dis_h_n net58 vgnd vcc_io sky130_fd_io__hvsbt_nand2
Xdm210 dm_h_n<2> and_dm01 dm_buf_dis vgnd vcc_io sky130_fd_io__hvsbt_nand2
Xdm10 dm_h_n<1> dm_h_n<0> nand_dm01 vgnd vcc_io sky130_fd_io__hvsbt_nand2
Xtripsel_nand net042 vtrip_sel_h tripsel_i_h_n vgnd vcc_io 
+ sky130_fd_io__hvsbt_nand2
.ENDS

.SUBCKT sky130_fd_io__com_inbuf_lv din out vgnd vpb vpwr
*.PININFO din:I vgnd:I vpb:I vpwr:I out:O
XI549 out din vgnd vgnd sky130_fd_pr__nfet_01v8 m=2 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI550 out din vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=3 w=5.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__com_inbuf_hv din out vcc_io vgnd
*.PININFO din:I vcc_io:I vgnd:I out:O
XI549 out din vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI550 out din vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__hvsbt_inv_x1_amux in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__or3_1 A B C X vgnd vnb vpb vpwr
*.PININFO A:I B:I C:I vgnd:I vnb:I vpb:I vpwr:I X:O
XMP0 vpwr A sndPA vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1 sndPA B sndPB vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP2 sndPB C y vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMIP3 X y vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN0 y A vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1 y B vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN2 y C vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMIN3 X y vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__nand3_1 A B C Y vgnd vnb vpb vpwr
*.PININFO A:I B:I C:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMP0 Y A vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1 Y B vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP2 Y C vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN0 Y A sndA vnb sky130_fd_pr__nfet_01v8 m=1 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1 sndA B sndB vnb sky130_fd_pr__nfet_01v8 m=1 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN2 sndB C vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amx_ls_bkp in in_b outb_hv pd_hv vgnd vhv
*.PININFO in:I in_b:I pd_hv:I vgnd:I vhv:I outb_hv:O
XI291 net54 net41 vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI287 net41 net54 vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI286 outb_hv net54 vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI283 net54 outb_hv vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI282 net41 outb_hv vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI278 net77 in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI276 outb_hv net54 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI273 net54 in_b vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI272 net41 outb_hv net77 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 net54 pd_hv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amx_inv2 A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XI73 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI72 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amx_inv4 A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XI75 Y A vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI74 Y A vda vda sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__inv_2 A Y vgnd vnb vpb vpwr
*.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMIN1 Y A vgnd vnb sky130_fd_pr__nfet_01v8 m=2 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMIP1 Y A vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=2 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amx_xor_lv A Ab B Bb out vgnd vnb vpb vpwr
*.PININFO A:I Ab:I B:I Bb:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI3 net39 B vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 out A net51 vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 net51 Bb vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out Ab net39 vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out A net64 vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 out Ab net76 vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI15 net76 Bb vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI14 net64 B vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amux_logic_decoder_lv amuxbusa_on amuxbusa_onb amuxbusb_on 
+ amuxbusb_onb analog_en analog_pol analog_sel out pd_on pd_onb pu_on pu_onb 
+ vccd vssd
*.PININFO analog_en:I analog_pol:I analog_sel:I out:I vccd:I vssd:I 
*.PININFO amuxbusa_on:O amuxbusa_onb:O amuxbusb_on:O amuxbusb_onb:O pd_on:O 
*.PININFO pd_onb:O pu_on:O pu_onb:O
XI357 amuxbusa_onb amuxbusa_on vssd vssd vccd vccd sky130_fd_io__inv_2
XI20 amuxbusb_onb amuxbusb_on vssd vssd vccd vccd sky130_fd_io__inv_2
XI16 out_b_i out_i vssd vssd vccd vccd sky130_fd_io__inv_2
XI348 out_i analog_pol_i pu_onb vssd vssd vccd vccd sky130_fd_io__nand2_1
XI19 analog_sel_i net56 amuxbusb_onb vssd vssd vccd vccd sky130_fd_io__nand2_1
XI26 out_b_i analog_pol_b pd_onb vssd vssd vccd vccd sky130_fd_io__nand2_1
XI18 net56 analog_sel_b amuxbusa_onb vssd vssd vccd vccd sky130_fd_io__nand2_1
XI17 out analog_en out_b_i vssd vssd vccd vccd sky130_fd_io__nand2_1
XI21 pd_onb pd_on vssd vssd vccd vccd sky130_fd_io__inv_1
XI31 analog_pol_b analog_pol_i vssd vssd vccd vccd sky130_fd_io__inv_1
XI28 analog_pol analog_pol_b vssd vssd vccd vccd sky130_fd_io__inv_1
XI32 analog_sel_b analog_sel_i vssd vssd vccd vccd sky130_fd_io__inv_1
XI22 pu_onb pu_on vssd vssd vccd vccd sky130_fd_io__inv_1
XI29 analog_sel analog_sel_b vssd vssd vccd vccd sky130_fd_io__inv_1
XI349 out_i out_b_i analog_pol_i analog_pol_b net56 vssd vssd vccd vccd 
+ sky130_fd_io__amx_xor_lv
.ENDS

.SUBCKT sky130_fd_io__amx_lslat_pd_1 in in_b out_vdda pd vccd vdda vssa
*.PININFO in:I in_b:I pd:I vccd:I vdda:I vssa:I out_vdda:O
XI11 latpu3 latpu4 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 latpu4 latpu3 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI59 out_vdda latpu3 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI21 latpu3 vccd net59 vssa sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI20 latpu4 vccd net55 vssa sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 latpu3 pd vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI167 out_vdda latpu3 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net59 in vssa vssa sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 net55 in_b vssa vssa sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amx_lslat in in_b out_vdda pd vccd vdda vssa
*.PININFO in:I in_b:I pd:I vccd:I vdda:I vssa:I out_vdda:O
XI11 latpu3 latpu4 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 latpu4 latpu3 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI59 out_vdda latpu3 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI21 latpu3 vccd net59 vssa sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI20 latpu4 vccd net55 vssa sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 latpu4 pd vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI167 out_vdda latpu3 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net59 in vssa vssa sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 net55 in_b vssa vssa sky130_fd_pr__nfet_01v8_lvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amx_ls_pdinv in in_b_pd in_pd pd_h vccd vccd_virt vssd
*.PININFO in:I pd_h:I vccd:I vccd_virt:I vssd:I in_b_pd:O in_pd:O
XI9 in_b_pd in vccd_virt vccd sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 in_pd in_b_pd vccd_virt vccd sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 in_pd pd_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 in_b_pd pd_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 in_pd in_b_pd vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 in_b_pd in vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amux_cntrl_logic_lv_sf analog_en analog_pol analog_sel 
+ ng_amx_vpmp_0 ng_amx_vpmp_1 ng_pad_vpmp_0 ng_pad_vpmp_1 nmid_vccd_0 
+ nmid_vccd_1 npd_vda out pd_vdda_n pd_vddio_n pg_amx_vda_0 pg_amx_vda_1 
+ pg_pad_vda_0 pg_pad_vda_1 ppu_vda vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I out:I pd_vdda_n:I pd_vddio_n:I 
*.PININFO vccd:I vdda:I vddio_q:I vssa:I vssd:I vswitch:I ng_amx_vpmp_0:O 
*.PININFO ng_amx_vpmp_1:O ng_pad_vpmp_0:O ng_pad_vpmp_1:O nmid_vccd_0:O 
*.PININFO nmid_vccd_1:O npd_vda:O pg_amx_vda_0:O pg_amx_vda_1:O pg_pad_vda_0:O 
*.PININFO pg_pad_vda_1:O ppu_vda:O
Xhld_i_h_inv1 pd_vdda_n pd_h_vdda vssa vdda sky130_fd_io__hvsbt_inv_x1_amux
XI515 pd_vddio_n pd_h_vddio vssd vddio_q sky130_fd_io__hvsbt_inv_x2
XI443 net234 net294 net178 vssd vssd vccd vccd sky130_fd_io__nand2_1
XI471 net228 net304 net171 vssd vssd vccd vccd sky130_fd_io__nand2_1
XI445 net178 amuxbusa_on nmid_vccd_0 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI436 net211 amuxbusa_onb net199 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI472 net171 amuxbusb_on nmid_vccd_1 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI473 net219 amuxbusb_onb net185 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI451 npd_vccd ppu_vccd_b nmid_vccd_1 net219 vssd vssd vccd vccd 
+ sky130_fd_io__or3_1
XI376 npd_vccd ppu_vccd_b nmid_vccd_0 net211 vssd vssd vccd vccd 
+ sky130_fd_io__or3_1
XI444 net178 switch_a_off vssd vssd vccd vccd sky130_fd_io__inv_1
XI448 net292 npd_vccd vssd vssd vccd vccd sky130_fd_io__inv_1
XI477 net171 switch_b_off vssd vssd vccd vccd sky130_fd_io__inv_1
XI449 net414 net234 vssd vssd vccd vccd sky130_fd_io__inv_1
XI476 net416 net228 vssd vssd vccd vccd sky130_fd_io__inv_1
XI392 switch_b_off switch_a_off pu_on net272 vssd vssd vccd vccd 
+ sky130_fd_io__nand3_1
XI435 switch_b_off switch_a_off pd_on net260 vssd vssd vccd vccd 
+ sky130_fd_io__nand3_1
XI381 net393 net394 net279 pd_h_vdda vssa vswitch sky130_fd_io__amx_ls_bkp
XI486 swtch_b_on swtch_b_off ng_pre_swtch_b pd_h_vdda vssa vswitch 
+ sky130_fd_io__amx_ls_bkp
XI447 npd_vda net292 vccd vssd sky130_fd_io__amx_inv2
XI496 ppu_vda ppu_vccd_b vccd vssd sky130_fd_io__amx_inv2
XI490 pg_amx_vda_1 net416 vccd vssd sky130_fd_io__amx_inv1
XI489 ng_amx_vpmp_1 net304 vccd vssd sky130_fd_io__amx_inv1
XI441 pg_amx_vda_0 net414 vccd vssd sky130_fd_io__amx_inv1
XI407 ng_amx_vpmp_0 net294 vccd vssd sky130_fd_io__amx_inv1
XI386 net363 pg_pad_vda_0 vdda vssa sky130_fd_io__amx_inv4
XI385 net363 pg_amx_vda_0 vdda vssa sky130_fd_io__amx_inv4
XI485 pg_pre_swtch_b pg_pad_vda_1 vdda vssa sky130_fd_io__amx_inv4
XI484 pg_pre_swtch_b pg_amx_vda_1 vdda vssa sky130_fd_io__amx_inv4
Xdecoder amuxbusa_on amuxbusa_onb amuxbusb_on amuxbusb_onb analog_en 
+ analog_pol analog_sel out pd_on pd_onb pu_on pu_onb vccd vssd 
+ sky130_fd_io__amux_logic_decoder_lv
XI439 net379 net380 pd_pre pd_h_vdda vccd_virt vswitch vssa 
+ sky130_fd_io__amx_lslat_pd_1
XI437 net393 net394 net363 pd_h_vdda vccd_virt vdda vssa sky130_fd_io__amx_lslat
XI497 net387 net386 net358 pd_h_vddio vccd_virt vddio_q vssd 
+ sky130_fd_io__amx_lslat
XI470 swtch_b_on swtch_b_off pg_pre_swtch_b pd_h_vdda vccd_virt vdda vssa 
+ sky130_fd_io__amx_lslat
XI498 net199 net394 net393 pd_h_vdda vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI500 net272 net387 net386 pd_h_vddio vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI501 net260 net380 net379 pd_h_vdda vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI499 net185 swtch_b_off swtch_b_on pd_h_vdda vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI502 vccd_virt pd_h_vdda vccd vccd sky130_fd_pr__pfet_g5v0d10v5 m=6 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI429 npd_vda pd_pre vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI431 ng_amx_vpmp_0 net279 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI517 npd_vda pd_pre vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI480 ng_amx_vpmp_1 ng_pre_swtch_b vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI479 ng_pad_vpmp_1 ng_pre_swtch_b vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI432 ng_pad_vpmp_0 net279 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI426 ppu_vda net358 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI415 ng_pad_vpmp_0 net279 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI519 npd_vda vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI428 ppu_vda net358 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI483 ng_pad_vpmp_1 ng_pre_swtch_b vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI482 ng_amx_vpmp_1 ng_pre_swtch_b vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI416 ng_amx_vpmp_0 net279 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI414 npd_vda pd_pre vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__amux_switch ag_hv ng_ag_vpmp ng_pad_vpmp nmid_vdda pad_hv_n0 
+ pad_hv_n1 pad_hv_n2 pad_hv_n3 pad_hv_p0 pad_hv_p1 pg_ag_vdda pg_pad_vdda 
+ vdda vddio_q vssa vssd
*.PININFO ng_ag_vpmp:I ng_pad_vpmp:I nmid_vdda:I pg_ag_vdda:I pg_pad_vdda:I 
*.PININFO vdda:I vddio_q:I vssa:I vssd:I ag_hv:B pad_hv_n0:B pad_hv_n1:B 
*.PININFO pad_hv_n2:B pad_hv_n3:B pad_hv_p0:B pad_hv_p1:B
XI56 vssa net109 sky130_fd_io__res75only_small
XI12 vssa net105 sky130_fd_io__res75only_small
XI26 ag_hv pg_ag_vdda mid vdda sky130_fd_pr__pfet_g5v0d10v5 m=4 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI22 pad_hv_p1 pg_pad_vdda mid vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI36 pad_hv_p0 pg_pad_vdda mid vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 ag_hv ng_ag_vpmp mid mid sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI35 pad_hv_n1 ng_pad_vpmp mid mid sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 pad_hv_n0 ng_pad_vpmp mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI57 mid_1 nmid_vdda net109 vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 mid nmid_vdda net105 vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI47 ag_hv ng_ag_vpmp mid_1 mid_1 sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI46 pad_hv_n3 ng_pad_vpmp mid_1 mid_1 sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI45 pad_hv_n2 ng_pad_vpmp mid_1 mid_1 sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_amux_sf amuxbus_a amuxbus_b analog_en analog_pol 
+ analog_sel out pad pd_vdda_n pd_vddio_n vccd vdda vddio_quiet vssa vssd 
+ vssio_quiet vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I out:I pd_vdda_n:I pd_vddio_n:I 
*.PININFO vccd:I vdda:I vddio_quiet:I vssa:I vssd:I vssio_quiet:I vswitch:I 
*.PININFO amuxbus_a:B amuxbus_b:B pad:B
XBBM_logic analog_en analog_pol analog_sel ng_amx_0 ng_amx_1 ng_pad_0 ng_pad_1 
+ nmid_0 nmid_1 pd_csd out pd_vdda_n pd_vddio_n pg_amx_0 pg_amx_1 pg_pad_0 
+ pg_pad_1 pu_csd vccd vdda vddio_quiet vssa vssd vswitch 
+ sky130_fd_io__amux_cntrl_logic_lv_sf
Xmux_a amuxbus_a ng_amx_0 ng_pad_0 nmid_0 net137 net137 net125 net125 net128 
+ net127 pg_amx_0 pg_pad_0 vdda vddio_quiet vssa vssd sky130_fd_io__amux_switch
Xmux_b amuxbus_b ng_amx_1 ng_pad_1 nmid_1 net137 net137 net125 net125 net128 
+ net127 pg_amx_1 pg_pad_1 vdda vddio_quiet vssa vssd sky130_fd_io__amux_switch
XI52 net148 pu_csd vddio_quiet vddio_quiet sky130_fd_pr__pfet_g5v0d10v5 m=3 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP_PU net152 pu_csd vddio_quiet vddio_quiet sky130_fd_pr__pfet_g5v0d10v5 m=4 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI49 net148 pd_csd vssio_quiet vssio_quiet sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN_PD net152 pd_csd vssio_quiet vssio_quiet sky130_fd_pr__nfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI26 net175 net137 sky130_fd_io__res75only_small
XI58 pad net127 sky130_fd_io__res75only_small
XI28 pad net128 sky130_fd_io__res75only_small
XI57 pad pad sky130_fd_io__res75only_small
XI27 net167 net125 sky130_fd_io__res75only_small
XI55 pad net175 sky130_fd_io__res75only_small
XI54 pad pad sky130_fd_io__res75only_small
XI53 pad net167 sky130_fd_io__res75only_small
XI40 pad net152 sky130_fd_io__res75only_small
XI39 pad net148 sky130_fd_io__res75only_small
.ENDS

.SUBCKT sky130_fd_io__com_ctl_ls_en hld_h_n hld_i_h in out_h rst_h_n vcc_io vpwr 
+ vssa vssd
*.PININFO hld_h_n:I hld_i_h:I in:I rst_h_n:I vcc_io:I vpwr:I vssa:I vssd:I 
*.PININFO out_h:O
XI34 in_i in_i_n vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 in_i_n in vpwr vpwr sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI70 fbk_n rst_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 in_i in_i_n vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out_h fbk_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI62 fbk hld_i_h vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 fbk_n hld_h_n net104 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI68 net104 in_i vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 in_i_n in vssd vssd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 fbk hld_h_n net84 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 fbk fbk_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI69 net84 in_i_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_ctl_lsbank analog_en analog_en_h dm<2> dm<1> dm<0> 
+ dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vdda_h hld_i_h 
+ hld_i_h_n inp_dis inp_dis_h inp_dis_h_n od_i_h vcc_io vdda vgnd vpwr vssa 
+ vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO analog_en:I dm<2>:I dm<1>:I dm<0>:I enable_vdda_h:I hld_i_h:I 
*.PININFO hld_i_h_n:I inp_dis:I od_i_h:I vcc_io:I vdda:I vgnd:I vpwr:I vssa:I 
*.PININFO vtrip_sel:I analog_en_h:O dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O 
*.PININFO dm_h_n<1>:O dm_h_n<0>:O inp_dis_h:O inp_dis_h_n:O vtrip_sel_h:O 
*.PININFO vtrip_sel_h_n:O
Xanalog_en_ls hld_i_h_n hld_i_h analog_en analog_en_h enable_vdda_h vdda vpwr 
+ vssa vgnd sky130_fd_io__com_ctl_ls_en
Xtrip_sel_st trip_sel_st_h od_i_h vgnd sky130_fd_io__tk_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h sky130_fd_io__tk_opti
Xdm_rst<2> dm_st_h<2> od_i_h vgnd sky130_fd_io__tk_opti
Xie_n_rst ie_n_rst_h vgnd od_i_h sky130_fd_io__tk_opti
Xdm_st<2> dm_rst_h<2> vgnd od_i_h sky130_fd_io__tk_opti
Xie_n_st ie_n_st_h od_i_h vgnd sky130_fd_io__tk_opti
Xdm_rst<1> dm_st_h<1> od_i_h vgnd sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> vgnd od_i_h sky130_fd_io__tk_opti
Xdm_st<1> dm_rst_h<1> vgnd od_i_h sky130_fd_io__tk_opti
XI337<1> dm_st_h<0> od_i_h vgnd sky130_fd_io__tk_opti
Xdm_ls<2> hld_i_h_n dm<2> dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> vcc_io vgnd 
+ vpwr sky130_fd_io__com_ctl_ls
Xdm_ls<1> hld_i_h_n dm<1> dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> vcc_io vgnd 
+ vpwr sky130_fd_io__com_ctl_ls
Xdm_ls<0> hld_i_h_n dm<0> dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> vcc_io vgnd 
+ vpwr sky130_fd_io__com_ctl_ls
Xinp_dis_ls hld_i_h_n inp_dis inp_dis_h inp_dis_h_n ie_n_rst_h ie_n_st_h 
+ vcc_io vgnd vpwr sky130_fd_io__com_ctl_ls
Xtrip_sel_ls hld_i_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n trip_sel_rst_h 
+ trip_sel_st_h vcc_io vgnd vpwr sky130_fd_io__com_ctl_ls
.ENDS

.SUBCKT sky130_fd_io__com_ctl_hld enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h 
+ hld_ovr od_i_h vcc_io vgnd vpwr
*.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h:O 
*.PININFO hld_i_h_n:O hld_i_ovr_h:O od_i_h:O
Xhld_ovr_ls net78 hld_ovr hld_ovr_h net46 vgnd vgnd vcc_io vgnd vpwr 
+ sky130_fd_io__com_ctl_ls
XI30 od_i_h hld_i_ovr_h_n hld_i_ovr_h vgnd vcc_io sky130_fd_io__hvsbt_nor
XI26 net78 hld_ovr_h hld_i_ovr_h_n vgnd vcc_io sky130_fd_io__hvsbt_nor
Xhld_i_h_inv4 net78 enable_vdda_h_n vgnd vcc_io sky130_fd_io__hvsbt_inv_x4
XI31 od_i_h_n od_i_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x4
Xhld_nand enable_h hld_h_n net73 vgnd vcc_io sky130_fd_io__hvsbt_nand2
Xod_h_inv enable_h od_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv1 net73 net78 vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
XI32 od_h od_i_h_n vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv8<1> enable_vdda_h_n hld_i_h_n_net<1> net018<0> net017<0> 
+ sky130_fd_io__hvsbt_inv_x8
Xhld_i_h_inv8<0> enable_vdda_h_n hld_i_h_n_net<0> net018<1> net017<1> 
+ sky130_fd_io__hvsbt_inv_x8
Rsky130_fd_pr__res_generic_m1<1> hld_i_h_n_net<1> hld_i_h_n sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
Rsky130_fd_pr__res_generic_m1<0> hld_i_h_n_net<0> hld_i_h_n sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
Rsky130_fd_pr__res_generic_m1_hld_i_h enable_vdda_h_n hld_i_h sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__gpio_ctl analog_en analog_en_h analog_en_vddio dm<2> dm<1> 
+ dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_h 
+ enable_inp_h enable_vdda_h hld_h_n hld_i_h_n hld_i_ovr_h hld_ovr inp_dis 
+ inp_dis_h_n inp_startup_en_h od_i_h vcc_io vdda vgnd vpwr vssa vtrip_sel 
+ vtrip_sel_h
*.PININFO analog_en:I dm<2>:I dm<1>:I dm<0>:I enable_h:I enable_inp_h:I 
*.PININFO enable_vdda_h:I hld_h_n:I hld_ovr:I inp_dis:I vcc_io:I vdda:I vgnd:I 
*.PININFO vpwr:I vssa:I vtrip_sel:I analog_en_h:O analog_en_vddio:O dm_h<2>:O 
*.PININFO dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O hld_i_h_n:O 
*.PININFO hld_i_ovr_h:O inp_dis_h_n:O inp_startup_en_h:O od_i_h:O vtrip_sel_h:O
XI56 od_i_h enable_inp_h net052 vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI51 analog_en_h enable_h net043 vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI57 net052 inp_startup_en_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
XI50 net043 analog_en_vddio vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xls_bank analog_en analog_en_h dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vdda_h hld_i_h hld_i_h_n inp_dis net49 
+ inp_dis_h_n od_i_h vcc_io vdda vgnd vpwr vssa vtrip_sel vtrip_sel_h net43 
+ sky130_fd_io__gpio_ctl_lsbank
Xhld_dis_blk enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr od_i_h 
+ vcc_io vgnd vpwr sky130_fd_io__com_ctl_hld
.ENDS

.SUBCKT sky130_fd_io__gpio_odrvr_sub force_hi_h_n force_lo_h force_lovol_h pad 
+ pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> 
+ tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io vssio_amx
*.PININFO force_hi_h_n:I force_lo_h:I force_lovol_h:I pd_h<3>:I pd_h<2>:I 
*.PININFO pd_h<1>:I pd_h<0>:I pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I 
*.PININFO vcc_io:I vgnd:I vgnd_io:I vssio_amx:I pad:O tie_hi_esd:B tie_lo_esd:B
Xpddrvr_strong force_lo_h force_lovol_h pad pd_h<3> pd_h<2> tie_lo_esd vcc_io 
+ vgnd_io vssio_amx sky130_fd_io__gpio_pddrvr_strong
Xpudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io vgnd 
+ sky130_fd_io__gpio_pudrvr_strong
Xpudrvr_weak weak_pad pu_h_n<0> vcc_io vgnd vcc_io sky130_fd_io__com_pudrvr_weak
Xpddrvr_weak weak_pad pd_h<0> vcc_io vgnd_io sky130_fd_io__gpio_pddrvr_weak
Xstrong_slow_pddrvr strong_slow_pad pd_h<1> vcc_io vgnd_io 
+ sky130_fd_io__gpio_pddrvr_strong_slow
Xstrong_slow_pudrvr strong_slow_pad pu_h_n<1> vcc_io vgnd vcc_io 
+ sky130_fd_io__com_pudrvr_strong_slow
Xres strong_slow_pad pad_r250 vgnd_io sky130_fd_io__com_res_strong_slow
Xres_weak weak_pad pad_r250 vgnd_io sky130_fd_io__com_res_weak
Xresd pad pad_r250 sky130_fd_io__res250only_small
.ENDS

.SUBCKT sky130_fd_io__gpio_odrvr force_hi_h_n force_lo_h force_lovol_h pad pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd 
+ tie_lo_esd vcc_io vgnd vgnd_io vssio_amx
*.PININFO force_hi_h_n:I force_lo_h:I force_lovol_h:I pd_h<3>:I pd_h<2>:I 
*.PININFO pd_h<1>:I pd_h<0>:I pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I 
*.PININFO vcc_io:I vgnd:I vgnd_io:I vssio_amx:I pad:O tie_hi_esd:O tie_lo_esd:O
Xbondpad pad vgnd_io sky130_fd_io__com_pad
Xodrvr force_hi_h_n force_lo_h force_lovol_h pad pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io 
+ vgnd vgnd_io vssio_amx sky130_fd_io__gpio_odrvr_sub
.ENDS

.SUBCKT sky130_fd_io__gpio_octl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n od_h pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h 
+ puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd vpwr vreg_en_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I od_h:I slow:I vcc_io:I vgnd:I vpwr:I vreg_en_h_n:I 
*.PININFO pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O puen_2or1_h:O puen_h<1>:O 
*.PININFO puen_h<0>:O slow_h:O slow_h_n:O
XI211 n<8> dm_h_n<1> puen_0_h vgnd vcc_io sky130_fd_io__hvsbt_nor
XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vcc_io sky130_fd_io__hvsbt_nor
XI210 dm_h<2> dm_h<0> n<8> vgnd vcc_io sky130_fd_io__hvsbt_xor
XI200 dm_h<2> dm_h<1> n<10> vgnd vcc_io sky130_fd_io__hvsbt_xor
XI185 dm_h_n<0> n<4> net119 vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI187 dm_h<1> dm_h<0> n<3> vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI203 n<10> dm_h<0> n<1> vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI204 n<9> dm_h_n<0> n<0> vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> puen_2or1_h vgnd vcc_io sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n puen_h<1> vgnd vcc_io sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n puen_h<0> vgnd vcc_io sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 pden_h_n<0> vgnd vcc_io sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 pden_h_n<1> vgnd vcc_io sky130_fd_io__hvsbt_inv_x2
XI377 puen_0_h puen_h0_n vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
XI374 net119 pden_h1 vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xls_slow hld_i_h_n slow slow_h slow_h_n od_h vgnd vcc_io vgnd vpwr 
+ sky130_fd_io__com_ctl_ls
.ENDS

.SUBCKT sky130_fd_io__com_opath_datoe drvhi_h drvlo_h_n hld_h_n hld_i_ovr_h od_h 
+ oe_h oe_n out vcc_io vgnd vpwr_ka
*.PININFO hld_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I vcc_io:I vgnd:I 
*.PININFO vpwr_ka:I drvhi_h:O drvlo_h_n:O oe_h:O
Xdat_ls hld_i_ovr_h out pd_dis_h pu_dis_h vgnd vgnd vcc_io vgnd vpwr_ka 
+ sky130_fd_io__gpio_dat_ls
Xoe_ls hld_i_ovr_h oe_n oe_h_n oe_h vgnd od_h vcc_io vgnd vpwr_ka 
+ sky130_fd_io__gpio_dat_ls
Xcclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io vgnd 
+ sky130_fd_io__com_cclat
.ENDS

.SUBCKT sky130_fd_io__gpio_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> en_fast_n<0> 
+ pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
Xmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin_fast<1> pd_h drvlo_h_n int_nor<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin_fast<0> pd_h drvlo_h_n int_nor<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI56 int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_pdpredrvr_strong drvlo_h_n pd_h<3> pd_h<2> pden_h_n 
+ slow_h vcc_io vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I slow_h:I vcc_io:I vgnd_io:I pd_h<3>:O 
*.PININFO pd_h<2>:O
XI77 en_fast2_n<1> pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI76 net76 pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> vcc_io sky130_fd_io__tk_opti
Xinv en_fast_h en_fast_h_n vgnd_io vcc_io sky130_fd_io__com_inv_x1_dnw
Xbias drvlo_h_n en_fast_h en_fast_h_n pbias_out pd_h<2> pden_h_n vcc_io 
+ vgnd_io sky130_fd_io__com_pdpredrvr_pbias
Xnor slow_h pden_h_n en_fast_h vgnd_io vcc_io sky130_fd_io__com_nor2_dnw
Xnr2 drvlo_h_n en_fast2_n<1> en_fast2_n<0> pd_h<3> pden_h_n vcc_io vgnd_io 
+ sky130_fd_io__gpio_pdpredrvr_strong_nr2
Xnr3 drvlo_h_n net76 net76 pd_h<2> pden_h_n vcc_io vgnd_io 
+ sky130_fd_io__gpio_pdpredrvr_strong_nr2
.ENDS

.SUBCKT sky130_fd_io__com_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XE1 net24 pu_h_n sky130_fd_io__tk_em1s
XRrespu1 int_res net24 sky130_fd_pr__res_generic_po m=1 w=0.33 l=11
XRrespu2 pu_h_n int_res sky130_fd_pr__res_generic_po m=1 w=0.33 l=4
Xmnin_fast<3> net24 drvhi_h int<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_fast<2> net24 drvhi_h int<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_fast<1> net24 drvhi_h int<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_fast<0> net24 drvhi_h int<0> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_slow1 n<2> puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_slow pu_h_n drvhi_h n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<3> int<3> en_fast<3> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<2> int<2> en_fast<2> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<1> int<1> en_fast<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h 
+ slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O
XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h sky130_fd_io__tk_opto
Xinv en_fast_h_n en_fast_h vgnd_io vcc_io sky130_fd_io__com_inv_x1_dnw
Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> 
+ pu_h_n<3> puen_h vcc_io vgnd_io sky130_fd_io__com_pupredrvr_strong_nd2
Xnd2a drvhi_h net54 net54 net54 net54 pu_h_n<2> puen_h vcc_io vgnd_io 
+ sky130_fd_io__com_pupredrvr_strong_nd2
Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io 
+ sky130_fd_io__com_pupredrvr_nbias
Xnand puen_h slow_h_n en_fast_h_n vgnd_io vcc_io sky130_fd_io__com_nand2_dnw
.ENDS

.SUBCKT sky130_fd_io__gpio_obpredrvr drvhi_h drvlo_h_n pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> 
+ puen_h<1> puen_h<0> slow_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I pden_h_n<1>:I pden_h_n<0>:I puen_h<1>:I 
*.PININFO puen_h<0>:I slow_h:I slow_h_n:I vcc_io:I vgnd_io:I pd_h<3>:O 
*.PININFO pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O 
*.PININFO pu_h_n<0>:O
Xpd_strong drvlo_h_n pd_h<3> pd_h<2> pden_h_n<1> slow_h vcc_io vgnd_io 
+ sky130_fd_io__gpio_pdpredrvr_strong
Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io 
+ sky130_fd_io__com_pupredrvr_weak
Xpd_weak drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io 
+ sky130_fd_io__com_pdpredrvr_weak
Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io 
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpd_strong_slow drvlo_h_n pd_h<1> pden_h_n<1> vcc_io vgnd_io 
+ sky130_fd_io__com_pdpredrvr_strong_slow
Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io 
+ sky130_fd_io__gpio_pupredrvr_strong
.ENDS

.SUBCKT sky130_fd_io__gpio_octl_dat dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h od_h oe_n out pd_h<3> pd_h<2> 
+ pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> slow slow_h_n vcc_io 
+ vgnd vgnd_io vpwr vpwr_ka
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I vpwr:I vpwr_ka:I drvhi_h:O pd_h<3>:O pd_h<2>:O pd_h<1>:O 
*.PININFO pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O slow_h_n:O
Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_h 
+ pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0> slow slow_h 
+ slow_h_n vcc_io vgnd vpwr vcc_io sky130_fd_io__gpio_octl
Xdatoe drvhi_h drvlo_h_n hld_i_h_n hld_i_ovr_h od_h oe_h oe_n out vcc_io vgnd 
+ vpwr_ka sky130_fd_io__com_opath_datoe
Xpredrvr drvhi_h drvlo_h_n pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> 
+ pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> 
+ slow_h slow_h_n vcc_io vgnd_io sky130_fd_io__gpio_obpredrvr
.ENDS

.SUBCKT sky130_fd_io__gpio_opath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hld_i_ovr_h od_h oe_n out pad slow tie_hi_esd tie_lo_esd 
+ vcc_io vgnd vgnd_io vpwr vpwr_ka vssio_amx
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I vpwr:I vpwr_ka:I vssio_amx:I pad:O tie_hi_esd:O 
*.PININFO tie_lo_esd:O
Xodrvr net68 net68 net68 pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io 
+ vssio_amx sky130_fd_io__gpio_odrvr
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n 
+ hld_i_ovr_h od_h oe_n out pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> slow slow_h_n vcc_io vgnd vgnd_io vpwr vpwr_ka 
+ sky130_fd_io__gpio_octl_dat
.ENDS

.SUBCKT sky130_fd_io__com_inbuf_ls en_h in_c in_t out_c out_t vgnd vpb vpwr
*.PININFO en_h:I in_c:I in_t:I vgnd:I vpb:I vpwr:I out_c:O out_t:O
XI534 out_t out_c vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_c out_t vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI536 out_c in_t vgnd_en vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_t in_c vgnd_en vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI552 vgnd_en en_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_inbuf_ls en_h en_h_n in_c in_t out_ls vgnd vpwr
*.PININFO en_h:I en_h_n:I in_c:I in_t:I vgnd:I vpwr:I out_ls:O
XI44 ls_out_n out_ls vgnd vgnd vpwr vpwr sky130_fd_io__gpio_inbuf_lvinv_x1
Xcom_ls en_h in_c in_t ls_out_n ls_out vgnd vpwr vpwr sky130_fd_io__com_inbuf_ls
XI561 ls_out_n en_h vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI54 ls_out en_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__com_ibuf_se en_h en_h_n ibufmux_out_h_n ibufmux_out_n in_h 
+ in_vt vcc_io vgnd vpwr_ka vtrip_sel_h_n
*.PININFO en_h:I en_h_n:I in_h:I in_vt:I vcc_io:I vgnd:I vpwr_ka:I 
*.PININFO vtrip_sel_h_n:I ibufmux_out_h_n:O ibufmux_out_n:O
Xhv_inv_1x out_h_wo_buf out_h_wo_buf_inv vcc_io vgnd vgnd 
+ sky130_fd_io__gpio_inbuf_hvinv_x1
Xhv_inv_4x<1> out_h_buf ibufmux_out_h_n net10<0> net12<0> net11<0> 
+ sky130_fd_io__gpio_inbuf_hvinv_x2
Xhv_inv_4x<0> out_h_buf ibufmux_out_h_n net10<1> net12<1> net11<1> 
+ sky130_fd_io__gpio_inbuf_hvinv_x2
Xhv_inv_2x out_h_wo_buf_inv out_h_buf vcc_io vgnd vgnd 
+ sky130_fd_io__gpio_inbuf_hvinv_x2
Xls en_h en_h_n out_h_n out_h_wo_buf out_ls vgnd vpwr_ka 
+ sky130_fd_io__gpio_inbuf_ls
Xlv_inv_x2 out_ls ibufmux_out_n vgnd vgnd vpwr_ka vpwr_ka 
+ sky130_fd_io__gpio_inbuf_lvinv_x2
Xbuf en_h in_h in_vt out_h_wo_buf out_h_n vcc_io vgnd vpwr_ka vtrip_sel_h_n 
+ sky130_fd_io__gpio_in_buf
.ENDS

.SUBCKT sky130_fd_io__gpio_ipath analog_en_h dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ inp_dis_h_n out out_h pad startup_en_h vcc_io vgnd vpwr_ka vtrip_sel_h
*.PININFO analog_en_h:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I inp_dis_h_n:I 
*.PININFO startup_en_h:I vcc_io:I vgnd:I vpwr_ka:I vtrip_sel_h:I out:O out_h:O 
*.PININFO pad:B
XLOGIC analog_en_h dm_h_n<2> dm_h_n<1> dm_h_n<0> inp_dis_h_n net37 net33 
+ startup_en_h tripsel_i_h tripsel_i_h_n vcc_io vgnd vtrip_sel_h 
+ sky130_fd_io__com_ictl_logic
Xesd pad in_h in_vt vcc_io vgnd tripsel_i_h sky130_fd_io__gpio_buf_localesd
Xibuf_se net33 net37 net51 net50 in_h in_vt vcc_io vgnd vpwr_ka tripsel_i_h_n 
+ sky130_fd_io__com_ibuf_se
Xmux_lv net50 out vgnd vpwr_ka vpwr_ka sky130_fd_io__com_inbuf_lv
Xmux_hv net51 out_h vcc_io vgnd sky130_fd_io__com_inbuf_hv
.ENDS

.SUBCKT sky130_fd_io__amux_cntrl_logic_lv analog_en analog_pol analog_sel 
+ ng_amx_vpmp_0 ng_amx_vpmp_1 ng_pad_vpmp_0 ng_pad_vpmp_1 nmid_vccd_0 
+ nmid_vccd_1 npd_vda out pd_vdda_n pd_vddio_n pg_amx_vda_0 pg_amx_vda_1 
+ pg_pad_vda_0 pg_pad_vda_1 ppu_vda vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I out:I pd_vdda_n:I pd_vddio_n:I 
*.PININFO vccd:I vdda:I vddio_q:I vssa:I vssd:I vswitch:I ng_amx_vpmp_0:O 
*.PININFO ng_amx_vpmp_1:O ng_pad_vpmp_0:O ng_pad_vpmp_1:O nmid_vccd_0:O 
*.PININFO nmid_vccd_1:O npd_vda:O pg_amx_vda_0:O pg_amx_vda_1:O pg_pad_vda_0:O 
*.PININFO pg_pad_vda_1:O ppu_vda:O
Xhld_i_h_inv1 pd_vdda_n pd_h_vdda vssa vdda sky130_fd_io__hvsbt_inv_x1_amux
XI515 pd_vddio_n pd_h_vddio vssd vddio_q sky130_fd_io__hvsbt_inv_x2
XI443 net228 net288 net172 vssd vssd vccd vccd sky130_fd_io__nand2_1
XI471 net222 net298 net165 vssd vssd vccd vccd sky130_fd_io__nand2_1
XI445 net172 amuxbusa_on nmid_vccd_0 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI436 net205 amuxbusa_onb net193 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI472 net165 amuxbusb_on nmid_vccd_1 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI473 net213 amuxbusb_onb net179 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI451 npd_vccd ppu_vccd_b nmid_vccd_1 net213 vssd vssd vccd vccd 
+ sky130_fd_io__or3_1
XI376 npd_vccd ppu_vccd_b nmid_vccd_0 net205 vssd vssd vccd vccd 
+ sky130_fd_io__or3_1
XI444 net172 switch_a_off vssd vssd vccd vccd sky130_fd_io__inv_1
XI448 net286 npd_vccd vssd vssd vccd vccd sky130_fd_io__inv_1
XI477 net165 switch_b_off vssd vssd vccd vccd sky130_fd_io__inv_1
XI449 net408 net228 vssd vssd vccd vccd sky130_fd_io__inv_1
XI476 net410 net222 vssd vssd vccd vccd sky130_fd_io__inv_1
XI392 switch_b_off switch_a_off pu_on net266 vssd vssd vccd vccd 
+ sky130_fd_io__nand3_1
XI435 switch_b_off switch_a_off pd_on net254 vssd vssd vccd vccd 
+ sky130_fd_io__nand3_1
XI381 net387 net388 net273 pd_h_vdda vssa vswitch sky130_fd_io__amx_ls_bkp
XI486 swtch_b_on swtch_b_off ng_pre_swtch_b pd_h_vdda vssa vswitch 
+ sky130_fd_io__amx_ls_bkp
XI447 npd_vda net286 vccd vssd sky130_fd_io__amx_inv2
XI496 ppu_vda ppu_vccd_b vccd vssd sky130_fd_io__amx_inv2
XI490 pg_amx_vda_1 net410 vccd vssd sky130_fd_io__amx_inv1
XI489 ng_amx_vpmp_1 net298 vccd vssd sky130_fd_io__amx_inv1
XI441 pg_amx_vda_0 net408 vccd vssd sky130_fd_io__amx_inv1
XI407 ng_amx_vpmp_0 net288 vccd vssd sky130_fd_io__amx_inv1
XI386 net357 pg_pad_vda_0 vdda vssa sky130_fd_io__amx_inv4
XI385 net357 pg_amx_vda_0 vdda vssa sky130_fd_io__amx_inv4
XI485 pg_pre_swtch_b pg_pad_vda_1 vdda vssa sky130_fd_io__amx_inv4
XI484 pg_pre_swtch_b pg_amx_vda_1 vdda vssa sky130_fd_io__amx_inv4
Xdecoder amuxbusa_on amuxbusa_onb amuxbusb_on amuxbusb_onb analog_en 
+ analog_pol analog_sel out pd_on pd_onb pu_on pu_onb vccd vssd 
+ sky130_fd_io__amux_logic_decoder_lv
XI439 net373 net374 pd_pre pd_h_vdda vccd_virt vswitch vssa 
+ sky130_fd_io__amx_lslat_pd_1
XI437 net387 net388 net357 pd_h_vdda vccd_virt vdda vssa sky130_fd_io__amx_lslat
XI497 net381 net380 net352 pd_h_vddio vccd_virt vddio_q vssd 
+ sky130_fd_io__amx_lslat
XI470 swtch_b_on swtch_b_off pg_pre_swtch_b pd_h_vdda vccd_virt vdda vssa 
+ sky130_fd_io__amx_lslat
XI498 net193 net388 net387 pd_h_vdda vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI500 net266 net381 net380 pd_h_vddio vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI501 net254 net374 net373 pd_h_vdda vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI499 net179 swtch_b_off swtch_b_on pd_h_vdda vccd vccd_virt vssd 
+ sky130_fd_io__amx_ls_pdinv
XI502 vccd_virt pd_h_vdda vccd vccd sky130_fd_pr__pfet_g5v0d10v5 m=6 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI429 npd_vda pd_pre vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI431 ng_amx_vpmp_0 net273 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI480 ng_amx_vpmp_1 ng_pre_swtch_b vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI479 ng_pad_vpmp_1 ng_pre_swtch_b vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI432 ng_pad_vpmp_0 net273 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI426 ppu_vda net352 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI415 ng_pad_vpmp_0 net273 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI428 ppu_vda net352 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI483 ng_pad_vpmp_1 ng_pre_swtch_b vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI482 ng_amx_vpmp_1 ng_pre_swtch_b vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI416 ng_amx_vpmp_0 net273 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI414 npd_vda pd_pre vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpio_amux amuxbus_a amuxbus_b analog_en analog_pol analog_sel 
+ out pad pd_vdda_n pd_vddio_n vccd vdda vddio_quiet vssa vssd vssio_quiet 
+ vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I out:I pd_vdda_n:I pd_vddio_n:I 
*.PININFO vccd:I vdda:I vddio_quiet:I vssa:I vssd:I vssio_quiet:I vswitch:I 
*.PININFO amuxbus_a:B amuxbus_b:B pad:B
XBBM_logic analog_en analog_pol analog_sel ng_amx_0 ng_amx_1 ng_pad_0 ng_pad_1 
+ nmid_0 nmid_1 pd_csd out pd_vdda_n pd_vddio_n pg_amx_0 pg_amx_1 pg_pad_0 
+ pg_pad_1 pu_csd vccd vdda vddio_quiet vssa vssd vswitch 
+ sky130_fd_io__amux_cntrl_logic_lv
Xmux_a amuxbus_a ng_amx_0 ng_pad_0 nmid_0 net212 net212 net200 net200 net203 
+ net202 pg_amx_0 pg_pad_0 vdda vddio_quiet vssa vssd sky130_fd_io__amux_switch
Xmux_b amuxbus_b ng_amx_1 ng_pad_1 nmid_1 net212 net212 net200 net200 net203 
+ net202 pg_amx_1 pg_pad_1 vdda vddio_quiet vssa vssd sky130_fd_io__amux_switch
XI52 net223 pu_csd vddio_quiet vddio_quiet sky130_fd_pr__pfet_g5v0d10v5 m=3 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP_PU net227 pu_csd vddio_quiet vddio_quiet sky130_fd_pr__pfet_g5v0d10v5 m=4 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI49 net223 pd_csd vssio_quiet vssio_quiet sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN_PD net227 pd_csd vssio_quiet vssio_quiet sky130_fd_pr__nfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI26 net250 net212 sky130_fd_io__res75only_small
XI58 pad net202 sky130_fd_io__res75only_small
XI28 pad net203 sky130_fd_io__res75only_small
XI57 pad pad sky130_fd_io__res75only_small
XI27 net242 net200 sky130_fd_io__res75only_small
XI55 pad net250 sky130_fd_io__res75only_small
XI54 pad pad sky130_fd_io__res75only_small
XI53 pad net242 sky130_fd_io__res75only_small
XI40 pad net227 sky130_fd_io__res75only_small
XI39 pad net223 sky130_fd_io__res75only_small
.ENDS

.SUBCKT sky130_fd_io__top_gpio amuxbus_a amuxbus_b analog_en analog_pol analog_sel 
+ dm<2> dm<1> dm<0> enable_h enable_inp_h enable_vdda_h hld_h_n hld_ovr in 
+ in_h inp_dis oe_n out pad pad_a_esd_0_h pad_a_esd_1_h pad_a_noesd_h slow 
+ tie_hi_esd tie_lo_esd vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q 
+ vswitch vtrip_sel
*.PININFO analog_en:I analog_pol:I analog_sel:I dm<2>:I dm<1>:I dm<0>:I 
*.PININFO enable_h:I enable_inp_h:I enable_vdda_h:I hld_h_n:I hld_ovr:I 
*.PININFO inp_dis:I oe_n:I out:I slow:I vtrip_sel:I in:O in_h:O tie_hi_esd:O 
*.PININFO tie_lo_esd:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_0_h:B 
*.PININFO pad_a_esd_1_h:B pad_a_noesd_h:B vccd:B vcchib:B vdda:B vddio:B 
*.PININFO vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xresd3 pad_a_esd_1_h net92 sky130_fd_io__res75only_small
Xresd1 net86 pad sky130_fd_io__res75only_small
Xresd4 net92 pad sky130_fd_io__res75only_small
Xresd2 pad_a_esd_0_h net86 sky130_fd_io__res75only_small
Xgpio_ctl analog_en analog_en_h analog_en_vddio dm<2> dm<1> dm<0> dm_h<2> 
+ dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_h enable_inp_h 
+ enable_vdda_h hld_h_n hld_i_h_n hld_i_ovr_h hld_ovr inp_dis inp_dis_h_n 
+ inp_startup_en_h od_i_h vddio_q vdda vssd vccd vssa vtrip_sel vtrip_sel_h 
+ sky130_fd_io__gpio_ctl
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_ovr_h od_i_h oe_n out pad slow tie_hi_esd tie_lo_esd vddio vssd vssio 
+ vccd vcchib vssa sky130_fd_io__gpio_opath
Xipath analog_en_h dm_h_n<2> dm_h_n<1> dm_h_n<0> inp_dis_h_n in in_h pad 
+ inp_startup_en_h vddio_q vssd vcchib vtrip_sel_h sky130_fd_io__gpio_ipath
Xamux amuxbus_a amuxbus_b analog_en analog_pol analog_sel out pad analog_en_h 
+ analog_en_vddio vccd vdda vddio_q vssa vssd vssio_q vswitch 
+ sky130_fd_io__gpio_amux
RS0<2> pad pad_a_noesd_h sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RS0<1> pad pad_a_noesd_h sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RS0<0> pad pad_a_noesd_h sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_hv_inv in out vddio_q vssd
*.PININFO in:I vddio_q:I vssd:I out:O
XI279 out in vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI277 out in vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_hv_nand2 in1 in2 out vddio_q vssd
*.PININFO in1:I in2:I vddio_q:I vssd:I out:O
XI280 out in2 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI279 out in1 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI277 out in1 net19 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI278 net19 in2 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_hv_nand3 in1 in2 in3 out vddio_q vssd
*.PININFO in1:I in2:I in3:I vddio_q:I vssd:I out:O
XI281 out in3 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI280 out in2 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI279 out in1 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI277 out in1 net27 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI282 net31 in3 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI278 net27 in2 net31 vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_hv_nor2 in1 in2 out vddio_q vssd
*.PININFO in1:I in2:I vddio_q:I vssd:I out:O
XI292 net10 in2 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI279 out in1 net10 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI277 out in1 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI293 out in2 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_decoder_5_32_cell in0 in1 in2 in3 in4 vddio_q 
+ vrefin vrefout vssd
*.PININFO in0:I in1:I in2:I in3:I in4:I vddio_q:I vrefin:I vssd:I vrefout:O
XI294 vrefin switch_en vrefout vssd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI283 vrefout net33 vrefin vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI280 switch_en net33 vddio_q vssd sky130_fd_io__gpiovrefv2_hv_inv
XI279 in3 in4 net37 vddio_q vssd sky130_fd_io__gpiovrefv2_hv_nand2
XI278 in0 in1 in2 net43 vddio_q vssd sky130_fd_io__gpiovrefv2_hv_nand3
XI277 net43 net37 switch_en vddio_q vssd sky130_fd_io__gpiovrefv2_hv_nor2
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_decoder_5_32 sel_h<4> sel_h<3> sel_h<2> sel_h<1> 
+ sel_h<0> selb_h<4> selb_h<3> selb_h<2> selb_h<1> selb_h<0> vddio_q vref<31> 
+ vref<30> vref<29> vref<28> vref<27> vref<26> vref<25> vref<24> vref<23> 
+ vref<22> vref<21> vref<20> vref<19> vref<18> vref<17> vref<16> vref<15> 
+ vref<14> vref<13> vref<12> vref<11> vref<10> vref<9> vref<8> vref<7> vref<6> 
+ vref<5> vref<4> vref<3> vref<2> vref<1> vref<0> vrefin vssd
*.PININFO sel_h<4>:I sel_h<3>:I sel_h<2>:I sel_h<1>:I sel_h<0>:I selb_h<4>:I 
*.PININFO selb_h<3>:I selb_h<2>:I selb_h<1>:I selb_h<0>:I vddio_q:I vref<31>:I 
*.PININFO vref<30>:I vref<29>:I vref<28>:I vref<27>:I vref<26>:I vref<25>:I 
*.PININFO vref<24>:I vref<23>:I vref<22>:I vref<21>:I vref<20>:I vref<19>:I 
*.PININFO vref<18>:I vref<17>:I vref<16>:I vref<15>:I vref<14>:I vref<13>:I 
*.PININFO vref<12>:I vref<11>:I vref<10>:I vref<9>:I vref<8>:I vref<7>:I 
*.PININFO vref<6>:I vref<5>:I vref<4>:I vref<3>:I vref<2>:I vref<1>:I 
*.PININFO vref<0>:I vssd:I vrefin:O
XI287 sel_h<0> selb_h<1> selb_h<2> selb_h<3> selb_h<4> vddio_q vref<1> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI277 selb_h<0> selb_h<1> selb_h<2> selb_h<3> selb_h<4> vddio_q vref<0> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI289 sel_h<0> sel_h<1> selb_h<2> selb_h<3> selb_h<4> vddio_q vref<3> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI288 selb_h<0> sel_h<1> selb_h<2> selb_h<3> selb_h<4> vddio_q vref<2> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI333 sel_h<0> selb_h<1> selb_h<2> sel_h<3> selb_h<4> vddio_q vref<9> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI332 selb_h<0> selb_h<1> selb_h<2> sel_h<3> selb_h<4> vddio_q vref<8> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI331 sel_h<0> sel_h<1> selb_h<2> sel_h<3> selb_h<4> vddio_q vref<11> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI330 selb_h<0> sel_h<1> selb_h<2> sel_h<3> selb_h<4> vddio_q vref<10> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI329 selb_h<0> sel_h<1> sel_h<2> sel_h<3> selb_h<4> vddio_q vref<14> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI328 sel_h<0> sel_h<1> sel_h<2> sel_h<3> selb_h<4> vddio_q vref<15> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI327 selb_h<0> selb_h<1> sel_h<2> sel_h<3> selb_h<4> vddio_q vref<12> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI349 selb_h<0> selb_h<1> sel_h<2> sel_h<3> sel_h<4> vddio_q vref<28> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI326 sel_h<0> selb_h<1> sel_h<2> sel_h<3> selb_h<4> vddio_q vref<13> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI321 selb_h<0> sel_h<1> sel_h<2> selb_h<3> selb_h<4> vddio_q vref<6> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI322 sel_h<0> sel_h<1> sel_h<2> selb_h<3> selb_h<4> vddio_q vref<7> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI323 selb_h<0> selb_h<1> sel_h<2> selb_h<3> selb_h<4> vddio_q vref<4> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI324 sel_h<0> selb_h<1> sel_h<2> selb_h<3> selb_h<4> vddio_q vref<5> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI358 sel_h<0> selb_h<1> selb_h<2> selb_h<3> sel_h<4> vddio_q vref<17> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI357 selb_h<0> selb_h<1> selb_h<2> selb_h<3> sel_h<4> vddio_q vref<16> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI356 sel_h<0> sel_h<1> selb_h<2> selb_h<3> sel_h<4> vddio_q vref<19> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI355 selb_h<0> sel_h<1> selb_h<2> selb_h<3> sel_h<4> vddio_q vref<18> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI354 selb_h<0> sel_h<1> sel_h<2> selb_h<3> sel_h<4> vddio_q vref<22> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI353 sel_h<0> sel_h<1> sel_h<2> selb_h<3> sel_h<4> vddio_q vref<23> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI352 selb_h<0> selb_h<1> sel_h<2> selb_h<3> sel_h<4> vddio_q vref<20> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI351 sel_h<0> selb_h<1> sel_h<2> selb_h<3> sel_h<4> vddio_q vref<21> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI350 sel_h<0> selb_h<1> sel_h<2> sel_h<3> sel_h<4> vddio_q vref<29> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI343 sel_h<0> selb_h<1> selb_h<2> sel_h<3> sel_h<4> vddio_q vref<25> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI344 selb_h<0> selb_h<1> selb_h<2> sel_h<3> sel_h<4> vddio_q vref<24> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI345 sel_h<0> sel_h<1> selb_h<2> sel_h<3> sel_h<4> vddio_q vref<27> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI346 selb_h<0> sel_h<1> selb_h<2> sel_h<3> sel_h<4> vddio_q vref<26> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI347 selb_h<0> sel_h<1> sel_h<2> sel_h<3> sel_h<4> vddio_q vref<30> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
XI348 sel_h<0> sel_h<1> sel_h<2> sel_h<3> sel_h<4> vddio_q vref<31> vrefin 
+ vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_res_ladder vddio_q vref<31> vref<30> vref<29> 
+ vref<28> vref<27> vref<26> vref<25> vref<24> vref<23> vref<22> vref<21> 
+ vref<20> vref<19> vref<18> vref<17> vref<16> vref<15> vref<14> vref<13> 
+ vref<12> vref<11> vref<10> vref<9> vref<8> vref<7> vref<6> vref<5> vref<4> 
+ vref<3> vref<2> vref<1> vref<0> vrefgen_en_h vrefgen_en_h_n vssd
*.PININFO vddio_q:I vrefgen_en_h:I vrefgen_en_h_n:I vssd:I vref<31>:O 
*.PININFO vref<30>:O vref<29>:O vref<28>:O vref<27>:O vref<26>:O vref<25>:O 
*.PININFO vref<24>:O vref<23>:O vref<22>:O vref<21>:O vref<20>:O vref<19>:O 
*.PININFO vref<18>:O vref<17>:O vref<16>:O vref<15>:O vref<14>:O vref<13>:O 
*.PININFO vref<12>:O vref<11>:O vref<10>:O vref<9>:O vref<8>:O vref<7>:O 
*.PININFO vref<6>:O vref<5>:O vref<4>:O vref<3>:O vref<2>:O vref<1>:O vref<0>:O
XI150 net81 vrefgen_en_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=10 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI191 net29 vrefgen_en_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=10 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI190 net99 vrefgen_en_h net29 vssd sky130_fd_pr__nfet_g5v0d10v5 m=10 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRI163 vref<26> vref<25> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI158 vref<28> vref<27> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI192 net99 net37 vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=2477.5
XRI209 vref<7> vref<8> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI162 vref<27> vref<26> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI197 vref<18> vref<19> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI160 vref<30> vref<29> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI161 vref<31> vref<30> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI196 vref<17> vref<18> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI213 vref<2> vref<3> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI198 vref<19> vref<20> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI157 net81 vref<31> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI215 vref<4> vref<5> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI199 vref<20> vref<21> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI201 vref<16> vref<15> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI212 vref<1> vref<2> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI195 vref<21> vref<22> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI193 vref<23> vref<24> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI194 vref<22> vref<23> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI207 vref<10> vref<9> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI164 vref<25> vref<24> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI204 vref<14> vref<13> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI205 vref<15> vref<14> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI206 vref<11> vref<10> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI159 vref<29> vref<28> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI200 vref<16> vref<17> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI214 vref<3> vref<4> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI378 net37 vref<0> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=2477.5
XRI216 vref<0> vref<1> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI210 vref<6> vref<7> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI211 vref<5> vref<6> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI202 vref<12> vref<11> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI208 vref<9> vref<8> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
XRI203 vref<13> vref<12> vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=350.09
.ENDS

.SUBCKT sky130_fd_io__gpiovrefv2_ctl enable_h hld_h_n sel<4> sel<3> sel<2> sel<1> 
+ sel<0> sel_h<4> sel_h<3> sel_h<2> sel_h<1> sel_h<0> selb_h<4> selb_h<3> 
+ selb_h<2> selb_h<1> selb_h<0> vccd vddio_q vrefgen_en vrefgen_en_h 
+ vrefgen_en_h_n vssd
*.PININFO enable_h:I hld_h_n:I sel<4>:I sel<3>:I sel<2>:I sel<1>:I sel<0>:I 
*.PININFO vccd:I vddio_q:I vrefgen_en:I vssd:I sel_h<4>:O sel_h<3>:O 
*.PININFO sel_h<2>:O sel_h<1>:O sel_h<0>:O selb_h<4>:O selb_h<3>:O selb_h<2>:O 
*.PININFO selb_h<1>:O selb_h<0>:O vrefgen_en_h:O vrefgen_en_h_n:O
Xhld_nand enable_h hld_h_n net32 vssd vddio_q sky130_fd_io__hvsbt_nand2
XI50 enable_h enable_h_n vssd vddio_q sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv1 net32 hld_i_h_n vssd vddio_q sky130_fd_io__hvsbt_inv_x1
XI353 hld_i_h_n vrefgen_en vrefgen_en_h vrefgen_en_h_n enable_h_n vssd vddio_q 
+ vssd vccd sky130_fd_io__com_ctl_ls
Xls<4> hld_i_h_n sel<4> sel_h<4> selb_h<4> enable_h_n vssd vddio_q vssd vccd 
+ sky130_fd_io__com_ctl_ls
Xls<3> hld_i_h_n sel<3> sel_h<3> selb_h<3> enable_h_n vssd vddio_q vssd vccd 
+ sky130_fd_io__com_ctl_ls
Xls<2> hld_i_h_n sel<2> sel_h<2> selb_h<2> enable_h_n vssd vddio_q vssd vccd 
+ sky130_fd_io__com_ctl_ls
Xls<1> hld_i_h_n sel<1> sel_h<1> selb_h<1> enable_h_n vssd vddio_q vssd vccd 
+ sky130_fd_io__com_ctl_ls
Xls<0> hld_i_h_n sel<0> sel_h<0> selb_h<0> enable_h_n vssd vddio_q vssd vccd 
+ sky130_fd_io__com_ctl_ls
.ENDS

.SUBCKT sky130_fd_io__top_gpiovrefv2 amuxbus_a amuxbus_b enable_h hld_h_n 
+ ref_sel<4> ref_sel<3> ref_sel<2> ref_sel<1> ref_sel<0> vccd vcchib vdda 
+ vddio vddio_q vinref vrefgen_en vssa vssd vssio vssio_q vswitch
*.PININFO enable_h:I hld_h_n:I ref_sel<4>:I ref_sel<3>:I ref_sel<2>:I 
*.PININFO ref_sel<1>:I ref_sel<0>:I vrefgen_en:I amuxbus_a:B amuxbus_b:B 
*.PININFO vccd:B vcchib:B vdda:B vddio:B vddio_q:B vinref:B vssa:B vssd:B 
*.PININFO vssio:B vssio_q:B vswitch:B
XI397 sel_h<4> sel_h<3> sel_h<2> sel_h<1> sel_h<0> selb_h<4> selb_h<3> 
+ selb_h<2> selb_h<1> selb_h<0> vddio_q vref<31> vref<30> vref<29> vref<28> 
+ vref<27> vref<26> vref<25> vref<24> vref<23> vref<22> vref<21> vref<20> 
+ vref<19> vref<18> vref<17> vref<16> vref<15> vref<14> vref<13> vref<12> 
+ vref<11> vref<10> vref<9> vref<8> vref<7> vref<6> vref<5> vref<4> vref<3> 
+ vref<2> vref<1> vref<0> vinref vssd sky130_fd_io__gpiovrefv2_decoder_5_32
XI276 vinref vrefgen_en_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI376 vddio_q vref<31> vref<30> vref<29> vref<28> vref<27> vref<26> vref<25> 
+ vref<24> vref<23> vref<22> vref<21> vref<20> vref<19> vref<18> vref<17> 
+ vref<16> vref<15> vref<14> vref<13> vref<12> vref<11> vref<10> vref<9> 
+ vref<8> vref<7> vref<6> vref<5> vref<4> vref<3> vref<2> vref<1> vref<0> 
+ vrefgen_en_h vrefgen_en_h_n vssd sky130_fd_io__gpiovrefv2_res_ladder
XI391 enable_h hld_h_n ref_sel<4> ref_sel<3> ref_sel<2> ref_sel<1> ref_sel<0> 
+ sel_h<4> sel_h<3> sel_h<2> sel_h<1> sel_h<0> selb_h<4> selb_h<3> selb_h<2> 
+ selb_h<1> selb_h<0> vccd vddio_q vrefgen_en vrefgen_en_h vrefgen_en_h_n vssd 
+ sky130_fd_io__gpiovrefv2_ctl
.ENDS

.SUBCKT sky130_fd_io__top_ground_padonlyv2 g_core g_pad
*.PININFO g_core:B g_pad:B
RI1 g_pad g_core sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__top_hvclamp drn_hvc ogc_hvc src_bdy_hvc
*.PININFO drn_hvc:B ogc_hvc:B src_bdy_hvc:B
Xpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc sky130_fd_pr__pfet_g5v0d10v5 m=50 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRrc_res g_pdpre net39 sky130_fd_pr__res_generic_po m=1 w=0.33 l=470
XRI38 net35 drn_hvc sky130_fd_pr__res_generic_po m=1 w=0.33 l=700
XRI37 net39 net35 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1550
Xclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=5.00 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=22 w=10.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__top_lvc_b2b bdy2_b2b drn_lvc1 drn_lvc2 ogc_lvc 
+ src_bdy_lvc1 src_bdy_lvc2 vssd
*.PININFO bdy2_b2b:B drn_lvc1:B drn_lvc2:B ogc_lvc:B src_bdy_lvc1:B 
*.PININFO src_bdy_lvc2:B vssd:B
XRI44 drn_lvc2 net66 sky130_fd_pr__res_generic_po m=1 w=0.33 l=900
XRI47 net66 net60 sky130_fd_pr__res_generic_po m=1 w=0.33 l=300
XRI46 g_pdpre_lvc2 net62 sky130_fd_pr__res_generic_po m=1 w=0.33 l=200
XRI45 net62 net60 sky130_fd_pr__res_generic_po m=1 w=0.33 l=720
XRrc_res g_pdpre_lvc1 drn_lvc1 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1950
Xncap src_bdy_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=15 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
Xpre_n1 g_nclamp_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=3 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI43 g_nclamp_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=2 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI58 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=6 w=5.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI60 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=1 w=5.00 
+ l=4.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI59 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=10 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
Xclamp_xtor drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=166 
+ w=7.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ area=0.063 perim=1.14
XI42 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=152 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI61 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 sky130_fd_pr__nfet_01v8 m=38 w=5.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI62 drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 sky130_fd_pr__nfet_01v8 m=20 w=5.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
Xpre_p1 g_nclamp_lvc1 g_pdpre_lvc1 drn_lvc1 drn_lvc1 sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI40 g_nclamp_lvc2 g_pdpre_lvc2 drn_lvc2 drn_lvc2 sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xesd bdy2_b2b src_bdy_lvc1 vssd sky130_fd_io__gnd2gnd_120x2_lv_isosub
.ENDS

.SUBCKT sky130_fd_io__top_lvclamp drn_lvc ogc_lvc src_bdy_lvc
*.PININFO drn_lvc:B ogc_lvc:B src_bdy_lvc:B
XRrc_res g_pdpre_lvc1 drn_lvc sky130_fd_pr__res_generic_po m=1 w=0.33 l=1950
Xncap src_bdy_lvc g_pdpre_lvc1 src_bdy_lvc src_bdy_lvc sky130_fd_pr__nfet_01v8 m=6 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
Xclamp_xtor drn_lvc g_nclamp_lvc1 src_bdy_lvc src_bdy_lvc sky130_fd_pr__nfet_01v8 m=204 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
Xpre_n1 g_nclamp_lvc1 g_pdpre_lvc1 src_bdy_lvc src_bdy_lvc sky130_fd_pr__nfet_01v8 m=2 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
XI57 src_bdy_lvc g_pdpre_lvc1 src_bdy_lvc src_bdy_lvc sky130_fd_pr__nfet_01v8 m=5 w=7.00 l=4.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpre_p1 g_nclamp_lvc1 g_pdpre_lvc1 drn_lvc drn_lvc sky130_fd_pr__pfet_01v8 m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__top_padv2 core pad
*.PININFO core:B pad:B
RI1 pad core sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__top_power_hvc_wpad amuxbus_a amuxbus_b drn_hvc ogc_hvc p_core 
+ p_pad src_bdy_hvc vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q 
+ vswitch
*.PININFO amuxbus_a:B amuxbus_b:B drn_hvc:B ogc_hvc:B p_core:B p_pad:B 
*.PININFO src_bdy_hvc:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B 
*.PININFO vssio:B vssio_q:B vswitch:B
Xpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc sky130_fd_pr__pfet_g5v0d10v5 m=50 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRrc_res g_pdpre net67 sky130_fd_pr__res_generic_po m=1 w=0.33 l=470
XRI38 net63 drn_hvc sky130_fd_pr__res_generic_po m=1 w=0.33 l=700
XRI37 net67 net63 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1550
Xclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=15 w=5.00 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc sky130_fd_pr__nfet_g5v0d10v5 m=22 w=10.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
RI13 p_pad p_core sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__top_power_padonlyv2 p_core p_pad
*.PININFO p_core:B p_pad:B
RI1 p_pad p_core sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__pwrdet_inv_4 A Y vgnd vnb vpb vpwr
*.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMIP1 Y A vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XMIN1 Y A vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__pwrdet_buf_4 A X vgnd vnb vpb vpwr
*.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I X:O
XMIN1 Ab A vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XMIN2 X Ab vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XMIP1 Ab A vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XMIP2 X Ab vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__pwrdet_lshv2hv_0 in out pd_hv vgnd vpwrin vpwrout
*.PININFO in:I pd_hv:I out:O vgnd:B vpwrin:B vpwrout:B
XI2 cross1 cross2 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 cross2 cross1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 net_158 pd_hvb vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 Ab in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI22 cross1 Ab net_158 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI21 cross2 Abb net_130 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 pd_hvb pd_hv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI16 net_138 cross2 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 cross1 pd_hv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 net_130 pd_hvb vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 Abb Ab vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 net120 cross1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 out net120 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 vgnd vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 Ab in vpwrin vpwrin sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI19 cross1 cross2 vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI15 net_138 cross2 vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 pd_hvb pd_hv vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 Abb Ab vpwrin vpwrin sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI18 cross2 cross1 vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 net120 cross1 vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 out net120 vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=8 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 vpwrout vpwrout vpwrout vpwrout sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__pwrdet_vddio out rst_por_hv_n vccd vddd vddio_q vssa vssd
*.PININFO rst_por_hv_n:I vccd:I vddd:I vddio_q:I vssa:I vssd:I out:O
XI7 net_1 out vssa vssa vddd vddd sky130_fd_io__pwrdet_inv_4
XI2 vddio_q net88 sky130_fd_io__res250only_small
XI21 pre_out out_1 net126 vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 vssa vddio_r vssa vssa sky130_fd_pr__nfet_05v0_nvt m=20 w=10.0 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI22 net126 rst_por_hv_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI16 net_1 out_1 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 net118 vddio_r net106 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 out_1 pre_out vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 vddio_b vddio_r net118 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 net106 vddio_r vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out_1 vddio_b vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI0 pre_out vddio_r vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI26 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI19 pre_out out_1 vddd vddd sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI15 vddd out_1 net_1 vddd sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI20 pre_out rst_por_hv_n vddd vddd sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI18 vccd vddio_r vddio_b vccd sky130_fd_pr__pfet_g5v0d10v5 m=8 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI14 out_1 pre_out vddd vddd sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 vddd vddd vddd vddd sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 vddd vddd vddd vddd sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XRI25 net88 vddio_r vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.3 l=278.07
.ENDS

.SUBCKT sky130_fd_io__pwrdet_vddd out vddd vddio_q vssa vssd
*.PININFO vddd:I vddio_q:I vssa:I out:O
XI0 vddd net100 sky130_fd_io__res250only_small
XI295 net194 n2 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI297 out net194 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI284 n2 n1 net117 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI285 n1 net129 p0 vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=4 w=7.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 net117 n1 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI20 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI19 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRI299 vssa vssa sky130_fd_pr__res_generic_po m=1 w=0.33 l=15.635
XRI2 p0 net138 vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.3 l=3150
XRI3 net132 vddio_q vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.3 l=1340
XRI12 vddd vddd vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.3 l=69.52
XRI9 net138 net132 sky130_fd_pr__res_generic_po m=1 w=0.33 l=1950
XRI11 net129 net100 vssd sky130_fd_pr__res_generic_nd__hv m=1 w=0.3 l=69.52
XI294 net194 n2 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI296 out net194 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI288 n2 n1 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=7.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI291 net182 net129 net178 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI292 net178 net129 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI289 n1 net129 net182 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 vssa net129 vssa vssa sky130_fd_pr__nfet_05v0_nvt m=15 w=10.0 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 vssa n2 vssa vssa sky130_fd_pr__nfet_05v0_nvt m=5 w=10.0 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI18 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI16 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI21 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI15 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI22 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__top_pwrdetv2 in1_vddd_hv in1_vddio_hv in2_vddd_hv 
+ in2_vddio_hv in3_vddd_hv in3_vddio_hv out1_vddd_hv out1_vddio_hv 
+ out2_vddd_hv out2_vddio_hv out3_vddd_hv out3_vddio_hv rst_por_hv_n 
+ tie_lo_esd vccd vddd1 vddd2 vddd_present_vddio_hv vddio_present_vddd_hv 
+ vddio_q vssa vssd vssio_q
*.PININFO in1_vddd_hv:I in1_vddio_hv:I in2_vddd_hv:I in2_vddio_hv:I 
*.PININFO in3_vddd_hv:I in3_vddio_hv:I rst_por_hv_n:I out1_vddd_hv:O 
*.PININFO out1_vddio_hv:O out2_vddd_hv:O out2_vddio_hv:O out3_vddd_hv:O 
*.PININFO out3_vddio_hv:O tie_lo_esd:O vddd_present_vddio_hv:O 
*.PININFO vddio_present_vddd_hv:O vccd:B vddd1:B vddd2:B vddio_q:B vssa:B 
*.PININFO vssd:B vssio_q:B
XI7 net166 net174 vssd vssd vddd1 vddd1 sky130_fd_io__pwrdet_inv_4
XI19 net178 net160 vssd vssd vddio_q vddio_q sky130_fd_io__pwrdet_inv_4
XI18 net178 vddd_present_vddio_hv vssd vssd vddio_q vddio_q 
+ sky130_fd_io__pwrdet_buf_4
XI2 net166 vddio_present_vddd_hv vssd vssd vddd1 vddd1 sky130_fd_io__pwrdet_buf_4
XI49 vssd tie_lo_esd sky130_fd_io__tk_tie_r_out_esd
XI17 in1_vddd_hv out1_vddio_hv net160 vssd vddd2 vddio_q 
+ sky130_fd_io__pwrdet_lshv2hv_0
XI16 in2_vddd_hv out2_vddio_hv net160 vssd vddd2 vddio_q 
+ sky130_fd_io__pwrdet_lshv2hv_0
XI3 in1_vddio_hv out1_vddd_hv net174 vssd vddio_q vddd1 
+ sky130_fd_io__pwrdet_lshv2hv_0
XI4 in2_vddio_hv out2_vddd_hv net174 vssd vddio_q vddd1 
+ sky130_fd_io__pwrdet_lshv2hv_0
XI5 in3_vddio_hv out3_vddd_hv net174 vssd vddio_q vddd1 
+ sky130_fd_io__pwrdet_lshv2hv_0
XI15 in3_vddd_hv out3_vddio_hv net160 vssd vddd2 vddio_q 
+ sky130_fd_io__pwrdet_lshv2hv_0
XI1 net166 rst_por_hv_n vccd vddd1 vddio_q vssa vssd sky130_fd_io__pwrdet_vddio
XI0 net178 vddd2 vddio_q vssa vssd sky130_fd_io__pwrdet_vddd
.ENDS

.SUBCKT sky130_fd_io__refgen_vdda_vswitch_ls in_h out_h out_h_n vddio_q vssa vswitch
*.PININFO in_h:I out_h:O out_h_n:O vddio_q:B vssa:B vswitch:B
XI446 in_i_h_n in_h vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 in_i_h in_i_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 out_h net66 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 out_h_n net58 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 net66 net58 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 net58 net66 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI449 in_i_h_n in_h vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI13 in_i_h in_i_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI17 out_h net66 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI25 out_h_n net58 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI0 net66 in_i_h vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 net58 in_i_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_ctl_vdda_ls_in_logic in in_dis out out_n vgnd vpb vpwr
*.PININFO in:I in_dis:I vgnd:I vpb:I vpwr:I out:O out_n:O
XI31 out in_dis vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 out_n in vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 out out_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 out_n in_dis vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI33 virt_pwr in_dis vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 virt_pwr in_dis vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 out_n in virt_pwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI34 out out_n virt_pwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_mux_and3 in_0 in_1 in_2 out vddio vssio
*.PININFO in_0:I in_1:I in_2:I out:O vddio:B vssio:B
XI31 net38 in_2 vssio vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 net34 in_0 net26 vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI34 out net34 vssio vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net26 in_1 net38 vssio sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 net34 in_2 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI35 out net34 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 net34 in_0 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 net34 in_1 vddio vddio sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_mux_dec sel<7> sel<6> sel<5> sel<4> sel<3> sel<2> 
+ sel<1> sel<0> vddio voh_sel_h<2> voh_sel_h<1> voh_sel_h<0> voh_sel_h_n<2> 
+ voh_sel_h_n<1> voh_sel_h_n<0> vssio
*.PININFO voh_sel_h<2>:I voh_sel_h<1>:I voh_sel_h<0>:I voh_sel_h_n<2>:I 
*.PININFO voh_sel_h_n<1>:I voh_sel_h_n<0>:I sel<7>:O sel<6>:O sel<5>:O 
*.PININFO sel<4>:O sel<3>:O sel<2>:O sel<1>:O sel<0>:O vddio:B vssio:B
XI12 voh_sel_h_n<2> voh_sel_h<1> voh_sel_h<0> sel<3> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI13 voh_sel_h<2> voh_sel_h_n<1> voh_sel_h<0> sel<5> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI16 voh_sel_h<2> voh_sel_h<1> voh_sel_h<0> sel<7> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI14 voh_sel_h<2> voh_sel_h_n<1> voh_sel_h_n<0> sel<4> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI15 voh_sel_h<2> voh_sel_h<1> voh_sel_h_n<0> sel<6> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI10 voh_sel_h_n<2> voh_sel_h_n<1> voh_sel_h<0> sel<1> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI11 voh_sel_h_n<2> voh_sel_h<1> voh_sel_h_n<0> sel<2> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
XI9 voh_sel_h_n<2> voh_sel_h_n<1> voh_sel_h_n<0> sel<0> vddio vssio 
+ sky130_fd_io__refgen_mux_and3
.ENDS

.SUBCKT sky130_fd_io__refgen_hvsbt_nand2 in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI3 out in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 out in1 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in1 net25 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net25 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_hvsbt_inv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_ctl_vdda_ls hld_h_n in in_n out_h out_h_n rst_h vdda 
+ vnb vpwr vssa
*.PININFO hld_h_n:I in:I in_n:I rst_h:I vdda:I vnb:I vpwr:I vssa:I out_h:O 
*.PININFO out_h_n:O
XI14 out_h_n fbk vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 out_h fbk_n vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 out_h_n fbk vssa vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out_h fbk_n vssa vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI58 net152 vpwr net0123 vnb sky130_fd_pr__nfet_05v0_nvt m=3 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnrst fbk rst_h vssa vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI59 net148 vpwr net0127 vnb sky130_fd_pr__nfet_05v0_nvt m=3 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 fbk_n hld_h_n net148 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 fbk hld_h_n net152 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk vssa vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 fbk fbk_n vssa vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 net0127 in vssa vnb sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 net0123 in_n vssa vnb sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_vddio_vswitch_ls in_i_h in_i_h_n out_h vssa vswitch
*.PININFO in_i_h:I in_i_h_n:I out_h:O vssa:B vswitch:B
XI16 out_h net67 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 net67 net59 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 net59 net67 vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 out_h net67 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI0 net67 in_i_h vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 net59 in_i_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_mux_and2 in_0 in_1 out vddio vssio
*.PININFO in_0:I in_1:I out:O vddio:B vssio:B
XI25 net20 out vssio vssio vddio vddio sky130_fd_io__refgen_hvsbt_inv_x1
XI24 in_1 in_0 net20 vssio vssio vddio vddio sky130_fd_io__refgen_hvsbt_nand2
.ENDS

.SUBCKT sky130_fd_io__refgen_ctl dft_refgen dft_refgen_vdda_n dft_refgen_vswitch 
+ enable_h enable_vdda_h hld_i_h_n hld_i_vpwr od_h sel_fb_mux<7> sel_fb_mux<6> 
+ sel_fb_mux<5> sel_fb_mux<4> sel_fb_mux<3> sel_fb_mux<2> sel_fb_mux<1> 
+ sel_fb_mux<0> sel_vdda_amuxbusa sel_vdda_amuxbusb sel_vdda_vref 
+ sel_vddio_amuxbusa sel_vddio_amuxbusb sel_vddio_vref vccd vdda vddio_q 
+ voh_sel<2> voh_sel<1> voh_sel<0> vref_sel<1> vref_sel<0> vref_sel_int vssa 
+ vssd vswitch
*.PININFO dft_refgen:I enable_h:I enable_vdda_h:I hld_i_h_n:I hld_i_vpwr:I 
*.PININFO voh_sel<2>:I voh_sel<1>:I voh_sel<0>:I vref_sel<1>:I vref_sel<0>:I 
*.PININFO dft_refgen_vdda_n:O dft_refgen_vswitch:O od_h:O sel_fb_mux<7>:O 
*.PININFO sel_fb_mux<6>:O sel_fb_mux<5>:O sel_fb_mux<4>:O sel_fb_mux<3>:O 
*.PININFO sel_fb_mux<2>:O sel_fb_mux<1>:O sel_fb_mux<0>:O sel_vdda_amuxbusa:O 
*.PININFO sel_vdda_amuxbusb:O sel_vdda_vref:O sel_vddio_amuxbusa:O 
*.PININFO sel_vddio_amuxbusb:O sel_vddio_vref:O vref_sel_int:O vccd:B vdda:B 
*.PININFO vddio_q:B vssa:B vssd:B vswitch:B
XI94 enable_vdda_h enable_vswitch_h net122 vdda vssa vswitch 
+ sky130_fd_io__refgen_vdda_vswitch_ls
XI53 vref_sel<0> hld_i_vpwr vref_sel0 vref_sel0_n vssd vccd vccd 
+ sky130_fd_io__refgen_ctl_vdda_ls_in_logic
XI50 vref_sel<1> hld_i_vpwr vref_sel1 vref_sel1_n vssd vccd vccd 
+ sky130_fd_io__refgen_ctl_vdda_ls_in_logic
XI54 dft_refgen hld_i_vpwr net151 net150 vssd vccd vccd 
+ sky130_fd_io__refgen_ctl_vdda_ls_in_logic
XI91 voh_sel<1> hld_i_vpwr voh_sel1 voh_sel1_n vssd vccd vccd 
+ sky130_fd_io__refgen_ctl_vdda_ls_in_logic
XI92 voh_sel<0> hld_i_vpwr voh_sel0 voh_sel0_n vssd vccd vccd 
+ sky130_fd_io__refgen_ctl_vdda_ls_in_logic
XI88 voh_sel<2> hld_i_vpwr voh_sel2 voh_sel2_n vssd vccd vccd 
+ sky130_fd_io__refgen_ctl_vdda_ls_in_logic
XI119 sel_fb_mux<7> sel_fb_mux<6> sel_fb_mux<5> sel_fb_mux<4> sel_fb_mux<3> 
+ sel_fb_mux<2> sel_fb_mux<1> sel_fb_mux<0> vswitch voh_sel_h<2> voh_sel_h<1> 
+ voh_sel_h<0> voh_sel_h_n<2> voh_sel_h_n<1> voh_sel_h_n<0> vssa 
+ sky130_fd_io__refgen_mux_dec
XI66 net209 enable_vdda_h sel_vdda_vref vssa vssa vdda vdda 
+ sky130_fd_io__refgen_hvsbt_nand2
XI67 net227 enable_vdda_h sel_vdda_amuxbusa vssa vssa vdda vdda 
+ sky130_fd_io__refgen_hvsbt_nand2
XI68 net233 enable_vdda_h sel_vdda_amuxbusb vssa vssa vdda vdda 
+ sky130_fd_io__refgen_hvsbt_nand2
XI52 vref_sel1_vdda vref_sel0_vdda net185 vssa vssa vdda vdda 
+ sky130_fd_io__refgen_hvsbt_nand2
XI51 vref_sel1_vdda vref_sel0_vdda_n net178 vssa vssa vdda vdda 
+ sky130_fd_io__refgen_hvsbt_nand2
XI22 net215 net239 vssa vssa vswitch vswitch sky130_fd_io__refgen_hvsbt_inv_x1
XI71 net185 net233 vssa vssa vdda vdda sky130_fd_io__refgen_hvsbt_inv_x1
XI70 net178 net227 vssa vssa vdda vdda sky130_fd_io__refgen_hvsbt_inv_x1
XI23 vref_sel1_vdda_n net221 vssa vssa vdda vdda sky130_fd_io__refgen_hvsbt_inv_x1
XI58 vref_sel1_vddio_n net215 vssa vssa vswitch vswitch 
+ sky130_fd_io__refgen_hvsbt_inv_x1
XI69 net221 net209 vssa vssa vdda vdda sky130_fd_io__refgen_hvsbt_inv_x1
XI436 vref_sel<1> vref_sel<0> net247 vssd vssd vccd vccd sky130_fd_io__nor2_1
XI444 net247 vref_sel_int vssd vssd vccd vccd sky130_fd_io__inv_1
XI13 hld_i_h_n_vswitch net151 net150 dft_refgen_vswitch net345 od_vswitch_h 
+ vswitch vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI38 hld_i_h_n_vdda net151 net150 net331 dft_refgen_vdda_n od_vdda_h vdda vssa 
+ vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI90 hld_i_h_n_vswitch voh_sel0 voh_sel0_n voh_sel_h<0> voh_sel_h_n<0> 
+ od_vswitch_h vswitch vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI49 hld_i_h_n_vdda vref_sel0 vref_sel0_n vref_sel0_vdda vref_sel0_vdda_n 
+ od_vdda_h vdda vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI48 hld_i_h_n_vdda vref_sel1 vref_sel1_n vref_sel1_vdda vref_sel1_vdda_n 
+ od_vdda_h vdda vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI21 hld_i_h_n_vswitch vref_sel1 vref_sel1_n vref_sel1_vddio vref_sel1_vddio_n 
+ od_vswitch_h vswitch vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI20 hld_i_h_n_vswitch vref_sel0 vref_sel0_n vref_sel0_vddio vref_sel0_vddio_n 
+ od_vswitch_h vswitch vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI57 hld_i_h_n_vswitch voh_sel1 voh_sel1_n voh_sel_h<1> voh_sel_h_n<1> 
+ od_vswitch_h vswitch vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI87 hld_i_h_n_vswitch voh_sel2 voh_sel2_n voh_sel_h<2> voh_sel_h_n<2> 
+ od_vswitch_h vswitch vssa vccd vssa sky130_fd_io__refgen_ctl_vdda_ls
XI105 net375 net371 vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104 net371 hld_i_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI96 od_vswitch_h enable_vswitch_h vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI242 od_h enable_h vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 od_vdda_h enable_vdda_h vdda vdda sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI107 net375 net371 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI106 net371 hld_i_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI241 od_h enable_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 od_vdda_h enable_vdda_h vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI97 od_vswitch_h enable_vswitch_h vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI61 net375 net371 net397 vssa vdda sky130_fd_io__refgen_vddio_vswitch_ls
XI59 net375 net371 net392 vssa vswitch sky130_fd_io__refgen_vddio_vswitch_ls
XI246 net397 enable_vdda_h hld_i_h_n_vdda vdda vssa sky130_fd_io__refgen_mux_and2
XI245 net392 enable_vswitch_h hld_i_h_n_vswitch vswitch vssa 
+ sky130_fd_io__refgen_mux_and2
XI63 enable_vswitch_h net239 sel_vddio_vref vswitch vssa 
+ sky130_fd_io__refgen_mux_and2
XI64 enable_vswitch_h net416 sel_vddio_amuxbusb vswitch vssa 
+ sky130_fd_io__refgen_mux_and2
XI24 enable_vswitch_h net421 sel_vddio_amuxbusa vswitch vssa 
+ sky130_fd_io__refgen_mux_and2
XI46 vref_sel0_vddio_n vref_sel1_vddio net421 vswitch vssa 
+ sky130_fd_io__refgen_mux_and2
XI47 vref_sel0_vddio vref_sel1_vddio net416 vswitch vssa 
+ sky130_fd_io__refgen_mux_and2
.ENDS

.SUBCKT sky130_fd_io__refgen_t_switch in out sel_vdda sel_vddio vdda vssa vswitch
*.PININFO in:I sel_vdda:I sel_vddio:I out:O vdda:B vssa:B vswitch:B
XI24 net056 sel_vdda_buf vssa vssa vdda vdda sky130_fd_io__refgen_hvsbt_inv_x1
XI114 sel_vdda net056 vssa vssa vdda vdda sky130_fd_io__refgen_hvsbt_inv_x1
XI28 sel_vddio net31 vssa vssa vswitch vswitch sky130_fd_io__refgen_hvsbt_inv_x1
XI27 net31 sel_vddio_buf vssa vssa vswitch vswitch 
+ sky130_fd_io__refgen_hvsbt_inv_x1
XI1 net26 sel_vdda in vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI21 out sel_vdda_buf net26 vdda sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 in sel_vddio net26 vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI22 net26 sel_vddio_buf out vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 net26 sel_vdda vssa vssa sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_dft dft_refgen_vdda_n dft_refgen_vswitch vdda vinref 
+ vinref_dft voutref voutref_dft vssa vswitch
*.PININFO dft_refgen_vdda_n:I dft_refgen_vswitch:I vinref:I voutref:I vdda:B 
*.PININFO vinref_dft:B voutref_dft:B vssa:B vswitch:B
XI229 voutref voutref_dft dft_refgen_vdda_n dft_refgen_vswitch vdda vssa 
+ vswitch sky130_fd_io__refgen_t_switch
XI228 vinref vinref_dft dft_refgen_vdda_n dft_refgen_vswitch vdda vssa vswitch 
+ sky130_fd_io__refgen_t_switch
.ENDS

.SUBCKT sky130_fd_io__refgen_com_ctl_ls hld_h_n in in_dis out_h out_h_n rst_h set_h 
+ vcc_io vgnd vpb vpwr
*.PININFO hld_h_n:I in:I in_dis:I rst_h:I set_h:I vcc_io:I vgnd:I vpb:I vpwr:I 
*.PININFO out_h:O out_h_n:O
XI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI34 in_i in_i_n virt_pwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 in_i_n in virt_pwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 virt_pwr in_dis vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI33 virt_pwr in_dis vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 in_i_n in_dis vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI58 net154 vpwr net114 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI59 net146 vpwr net118 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 fbk_n hld_h_n net146 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 in_i in_dis vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 fbk hld_h_n net154 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 net118 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 net114 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_vpwrka_ls in_h in_h_n out_n vgnd vpwr_ka
*.PININFO in_h:I in_h_n:I vgnd:I vpwr_ka:I out_n:O
XI4 out_n net30 vgnd vgnd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI334 net30 in_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 net35 in_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI187 out_n net30 vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 net35 net30 vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 net30 net35 vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_em1s a b
*.PININFO a:B b:B
RI1 a net8 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI2 b net8 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__refgen_em1o a b
*.PININFO a:B b:B
RI1 a net11 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI2 b net7 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__refgen_opti out spd spu
*.PININFO out:B spd:B spu:B
Xe1 out spu sky130_fd_io__refgen_em1s
Xe2 spd out sky130_fd_io__refgen_em1o
.ENDS

.SUBCKT sky130_fd_io__refgen_inv_x8 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=8 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=8 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_inv_x4 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_inv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_nand2 in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI3 out in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 out in1 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in1 net25 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net25 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__inv_p in0 out vgnd vnb vpb vpwr
*.PININFO in0:I vgnd:I vnb:I vpb:I vpwr:I out:O
X8 out in0 vgnd vnb sky130_fd_pr__nfet_01v8 m=nm w=nw l=nl mult=1 sa=nsa sb=nsb sd=nsd 
+ topography=normal area=0.063 perim=1.14
X7 out in0 vpwr vpb sky130_fd_pr__pfet_01v8 m=pm w=pw l=pl mult=1 sa=psa sb=psb sd=psd 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_in_ctl_ls_out in_c in_t out_c out_t vgnd vpb vpwr
*.PININFO in_c:I in_t:I vgnd:I vpb:I vpwr:I out_c:O out_t:O
XI35 out_c_n out_c vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 psa=265e-3 
+ pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 nw=1.00 nm=1
XI36 out_t_n out_t vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 psa=265e-3 
+ pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 nw=1.00 nm=1
XI536 out_t_n in_t vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_c_n in_c vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI534 out_c_n out_t_n vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_t_n out_c_n vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_lvlp_inv_x4 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI1 out in vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=4 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 out in vgnd vnb sky130_fd_pr__nfet_01v8 m=4 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_ctl_hld hld_h_n hld_i_h_n hld_i_vpwr od_h vcc_io vgnd 
+ vpb vpwr
*.PININFO hld_h_n:I od_h:I vcc_io:I vgnd:I vpb:I vpwr:I hld_i_h_n:O 
*.PININFO hld_i_vpwr:O
Xhld_i_h_inv8<1> hld_i_h hld_i_h_n vgnd vgnd vcc_io vcc_io
+ sky130_fd_io__refgen_inv_x8
Xhld_i_h_inv8<0> hld_i_h hld_i_h_n vgnd vgnd vcc_io vcc_io
+ sky130_fd_io__refgen_inv_x8
Xhld_i_h_inv4 hld_i_h_n_ls hld_i_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_inv_x4
Xod_h_inv od_h od_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x1
Xhld_i_h_inv1 hld_i_h_ls hld_i_h_n_ls vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_inv_x1
Xhld_nand od_h_n hld_h_n hld_i_h_ls vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
Xhld_i_vpwr_ls hld_i_h_n_ls hld_i_h_ls hld_i_vpwr_n net24 vgnd vpb vpwr 
+ sky130_fd_io__refgen_in_ctl_ls_out
Xhld_i_vpwr_inv hld_i_vpwr_n hld_i_vpwr vgnd vgnd vpb vpwr 
+ sky130_fd_io__refgen_lvlp_inv_x4
.ENDS

.SUBCKT sky130_fd_io__refgen_in_xlators biasen_n hld_h_n hld_i_h_n hld_i_vpwr 
+ ibuf_sel ibuf_sel_h ibuf_sel_h_n ls_in_h ls_in_h_n od_h vcc_a vcc_io vgnd 
+ vpb vpwr vpwr_ka vref_sel vref_sel_h vref_sel_h_n vreg_en vreg_en_h 
+ vreg_en_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO hld_h_n:I ibuf_sel:I ls_in_h:I ls_in_h_n:I od_h:I vref_sel:I 
*.PININFO vreg_en:I vtrip_sel:I biasen_n:O hld_i_h_n:O hld_i_vpwr:O 
*.PININFO ibuf_sel_h:O ibuf_sel_h_n:O vref_sel_h:O vref_sel_h_n:O vreg_en_h:O 
*.PININFO vreg_en_h_n:O vtrip_sel_h:O vtrip_sel_h_n:O vcc_a:B vcc_io:B vgnd:B 
*.PININFO vpb:B vpwr:B vpwr_ka:B
Xls_vref_sel hld_i_h_n vref_sel hld_i_vpwr vref_sel_h vref_sel_h_n 
+ ref_sel_rst_h ref_sel_st_h vcc_a vgnd vpb vpwr sky130_fd_io__refgen_com_ctl_ls
Xls_vtrip_sel hld_i_h_n vtrip_sel hld_i_vpwr vtrip_sel_h vtrip_sel_h_n 
+ trip_sel_rst_h trip_sel_st_h vcc_a vgnd vpb vpwr sky130_fd_io__refgen_com_ctl_ls
Xls_vreg_en hld_i_h_n vreg_en hld_i_vpwr vreg_en_h vreg_en_h_n net86 net89 
+ vcc_a vgnd vpb vpwr sky130_fd_io__refgen_com_ctl_ls
Xls_ibuf_sel hld_i_h_n ibuf_sel hld_i_vpwr ibuf_sel_h ibuf_sel_h_n 
+ buf_sel_rst_h buf_sel_st_h vcc_a vgnd vpb vpwr sky130_fd_io__refgen_com_ctl_ls
Xls_vreg_en_ka ls_in_h ls_in_h_n biasen_n vgnd vpwr_ka 
+ sky130_fd_io__refgen_vpwrka_ls
XI458 ref_sel_st_h od_h vgnd sky130_fd_io__refgen_opti
XI459 ref_sel_rst_h vgnd od_h sky130_fd_io__refgen_opti
XI471 net89 od_h vgnd sky130_fd_io__refgen_opti
XI470 net86 vgnd od_h sky130_fd_io__refgen_opti
Xbuf_sel_rst buf_sel_rst_h vgnd od_h sky130_fd_io__refgen_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_h sky130_fd_io__refgen_opti
Xbuf_sel_st buf_sel_st_h od_h vgnd sky130_fd_io__refgen_opti
Xtrip_sel_st trip_sel_st_h od_h vgnd sky130_fd_io__refgen_opti
Xhld_blk hld_h_n hld_i_h_n hld_i_vpwr od_h vcc_io vgnd vpb vpwr 
+ sky130_fd_io__refgen_ctl_hld
.ENDS

.SUBCKT sky130_fd_io__refgen_opamp_stage_1_res b r1 r2 vgnd
*.PININFO vgnd:I b:B r1:B r2:B
XRI345 net61 net62 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI1 net58 net61 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI2 net55 net58 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI3 r1 net49 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI4 net49 net55 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI5 net46 net40 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI6 net43 net46 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI7 net40 net37 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI8 net37 net34 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI9 net34 net62 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI10 net31 net5 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI11 net28 net31 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI12 net25 net28 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI13 r2 net19 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI14 net19 net25 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI15 net16 net10 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI16 net43 net16 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI17 net10 net7 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI18 net7 net4 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI19 net4 net5 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI36 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI35 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI34 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI33 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI32 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI37 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI38 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI39 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI40 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
XRI41 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.675
.ENDS

.SUBCKT sky130_fd_io__refgen_opamp_stage_1 en_inpop_h ibuf_sel_h_n inn inp ngate 
+ out vcc vgnd
*.PININFO en_inpop_h:I ibuf_sel_h_n:I inn:I inp:I vcc:I vgnd:I out:O ngate:B
XI345 vgnd out net186 vgnd sky130_fd_io__refgen_opamp_stage_1_res
XI153 net130 vsource sky130_fd_io__refgen_em1o
XI220 net150 vsource sky130_fd_io__refgen_em1o
XI223 net142 vsource sky130_fd_io__refgen_em1o
XI214 net126 net111 sky130_fd_io__refgen_em1o
XI211 net126 net77 sky130_fd_io__refgen_em1o
XI250 vgnd net167 sky130_fd_io__refgen_em1o
XI255 net171 out sky130_fd_io__refgen_em1o
XI253 net163 out sky130_fd_io__refgen_em1o
XI252 net163 vgnd sky130_fd_io__refgen_em1s
XI215 vcc net111 sky130_fd_io__refgen_em1s
XI212 vcc net77 sky130_fd_io__refgen_em1s
XI228 net195 net138 sky130_fd_io__refgen_em1s
XE3 net195 net134 sky130_fd_io__refgen_em1s
XI467 out net186 sky130_fd_io__refgen_em1s
XI254 net171 vgnd sky130_fd_io__refgen_em1s
XI243 out net167 sky130_fd_io__refgen_em1s
XMP<1> net186 net77 vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<2> net126 net126 vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<0> net126 net111 vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<3> net186 net126 vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI217<3> net126 en_inpop_h vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI216<3> vcc vcc vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI230<3> net142 ngate net138 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> vsource ngate net195 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<2> net150 ngate net195 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> net130 ngate net195 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<3> net142 ngate net195 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI227 net138 en_inpop_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI224 net134 en_inpop_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI229<1> net130 ngate net134 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI219 net186 vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN2 net186 inn vsource vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1 net126 inp vsource vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI218 net126 vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI232 net186 ibuf_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI256 vgnd net171 vgnd vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI209 vgnd net167 vgnd vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI241 vgnd net163 vgnd vgnd sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_c r0 r1 vnb
*.PININFO r0:B r1:B vnb:B
XI315 net49 net46 sky130_fd_io__refgen_em1o
XI314 net52 net49 sky130_fd_io__refgen_em1o
XI313 r1 net52 sky130_fd_io__refgen_em1o
XI312 net55 net43 sky130_fd_io__refgen_em1o
XI311 net43 net37 sky130_fd_io__refgen_em1o
XI467 net37 r0 sky130_fd_io__refgen_em1o
XRI316 net40 net55 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<13> r1 net52 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<12> net52 net49 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<11> net49 net46 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<4> net55 net43 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI317<1> net46 net40 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<1> net43 net37 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<0> net37 r0 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_d r0 r1 vnb
*.PININFO r0:B r1:B vnb:B
XI315 net49 net46 sky130_fd_io__refgen_em1o
XI314 net52 net49 sky130_fd_io__refgen_em1o
XI313 r1 net52 sky130_fd_io__refgen_em1o
XI312 net55 net43 sky130_fd_io__refgen_em1o
XI311 net43 net37 sky130_fd_io__refgen_em1o
XI467 net37 r0 sky130_fd_io__refgen_em1o
XRI316 net40 net55 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<13> r1 net52 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<12> net52 net49 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<11> net49 net46 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<4> net55 net43 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI317<1> net46 net40 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<1> net43 net37 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR<0> net37 r0 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_g r0 r1 vnb
*.PININFO r0:B r1:B vnb:B
XI320 net41 net53 sky130_fd_io__refgen_em1o
XI319 net53 r0 sky130_fd_io__refgen_em1o
XI325 net62 net59 sky130_fd_io__refgen_em1o
XI324 net65 net62 sky130_fd_io__refgen_em1o
XI323 r1 net65 sky130_fd_io__refgen_em1o
XI467 net44 net41 sky130_fd_io__refgen_em1o
XRR1<0> net53 r0 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<5> net47 net77 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<9> net73 net74 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<8> net74 net71 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<10> net59 net73 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.955
XRR1<13> r1 net65 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<12> net65 net62 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<11> net62 net59 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<7> net71 net56 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<1> net41 net53 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<4> net77 net50 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<6> net56 net47 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<3> net50 net44 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<2> net44 net41 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_h r0 r1 vnb
*.PININFO r0:B r1:B vnb:B
XI320 net41 net53 sky130_fd_io__refgen_em1o
XI319 net53 r0 sky130_fd_io__refgen_em1o
XI325 net62 net59 sky130_fd_io__refgen_em1o
XI324 net65 net62 sky130_fd_io__refgen_em1o
XI323 r1 net65 sky130_fd_io__refgen_em1o
XI467 net44 net41 sky130_fd_io__refgen_em1o
XRR1<0> net53 r0 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<5> net47 net77 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<9> net73 net74 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<8> net74 net71 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<10> net59 net73 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.955
XRR1<13> r1 net65 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<12> net65 net62 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<11> net62 net59 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<7> net71 net56 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<1> net41 net53 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<4> net77 net50 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<6> net56 net47 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<3> net50 net44 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<2> net44 net41 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_i r0 r1 vnb
*.PININFO r0:B r1:B vnb:B
XI320 net41 net53 sky130_fd_io__refgen_em1o
XI319 net53 r0 sky130_fd_io__refgen_em1o
XI325 net62 net59 sky130_fd_io__refgen_em1o
XI324 net65 net62 sky130_fd_io__refgen_em1o
XI323 r1 net65 sky130_fd_io__refgen_em1o
XI467 net44 net41 sky130_fd_io__refgen_em1o
XRR1<0> net53 r0 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<5> net47 net77 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<9> net73 net74 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<8> net74 net71 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<10> net59 net73 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.955
XRR1<13> r1 net65 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<12> net65 net62 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<11> net62 net59 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<7> net71 net56 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<1> net41 net53 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<4> net77 net50 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<6> net56 net47 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<3> net50 net44 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRR1<2> net44 net41 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
.ENDS

.SUBCKT sky130_fd_io__refgen_in_lpf ibuf_sel_h_n in out vcc_a vgnd
*.PININFO ibuf_sel_h_n:I in:I vcc_a:I vgnd:I out:O
XI102 vcc_a net73 sky130_fd_io__refgen_em1s
XI118 net126 net114 sky130_fd_io__refgen_em1s
XI119 vcc_a net63 sky130_fd_io__refgen_em1s
XI120 vcc_a net75 sky130_fd_io__refgen_em1s
XI44 net87 out sky130_fd_io__refgen_em1s
XI101 net100 out sky130_fd_io__refgen_em1s
XI117 net114 out sky130_fd_io__refgen_em1s
XI77 net118 net100 sky130_fd_io__refgen_em1s
XI76 vcc_a net57 sky130_fd_io__refgen_em1s
XI572 net135 out sky130_fd_io__refgen_em1o
XI16 net97 in sky130_fd_io__refgen_em1o
XI17 net95 net97 sky130_fd_io__refgen_em1o
XI114 net75 net126 sky130_fd_io__refgen_em1o
XI18 net91 net95 sky130_fd_io__refgen_em1o
XI19 net89 net91 sky130_fd_io__refgen_em1o
XI20 net87 net89 sky130_fd_io__refgen_em1o
XI21 net85 net87 sky130_fd_io__refgen_em1o
XI22 net83 net85 sky130_fd_io__refgen_em1o
XI23 net81 net83 sky130_fd_io__refgen_em1o
XI24 net79 net81 sky130_fd_io__refgen_em1o
XI25 net77 net79 sky130_fd_io__refgen_em1o
XI116 net75 vgnd sky130_fd_io__refgen_em1o
XI99 net73 net100 sky130_fd_io__refgen_em1o
XI46 net79 out sky130_fd_io__refgen_em1o
XI45 net83 out sky130_fd_io__refgen_em1o
XI43 net91 out sky130_fd_io__refgen_em1o
XI42 net97 out sky130_fd_io__refgen_em1o
XI115 net63 net114 sky130_fd_io__refgen_em1o
XI113 net63 vgnd sky130_fd_io__refgen_em1o
XI100 net73 vgnd sky130_fd_io__refgen_em1o
XI79 net57 vgnd sky130_fd_io__refgen_em1o
XI78 net57 net118 sky130_fd_io__refgen_em1o
XI571 net135 ibuf_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI90 net114 net63 net114 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI89 net126 net75 net126 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI80 net100 net73 net100 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI75 net118 net57 net118 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRI15 net79 net77 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI14 net81 net79 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI13 net83 net81 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI12 net85 net83 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI11 net87 net85 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI10 net87 net89 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI9 net89 net91 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI8 net91 net95 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI7 net95 net97 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI6 net97 in vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
.ENDS

.SUBCKT sky130_fd_io__refgen_ls in in_n out vcc_io vgnd
*.PININFO in:I in_n:I vcc_io:I vgnd:I out:O
XI45 out out_t_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI536 out_t_n in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 net37 in_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI534 net37 out_t_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_t_n net37 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI44 out out_t_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_vinref_1 ibuf_sel_h ibuf_sel_h_n in_lpf 
+ sel_vcc_io sel_vcc_io_0p4 vcc_a vcc_io vcc_io_0p5 vgnd vinref
*.PININFO ibuf_sel_h:I ibuf_sel_h_n:I in_lpf:I sel_vcc_io:I sel_vcc_io_0p4:I 
*.PININFO vgnd:I vinref:O vcc_a:B vcc_io:B vcc_io_0p5:B
XR<1> net75 net78 vgnd sky130_fd_io__refgen_res_ntwk_c
XR<0> net76 net75 vgnd sky130_fd_io__refgen_res_ntwk_c
XR<2> net78 net72 vgnd sky130_fd_io__refgen_res_ntwk_c
XR<3> net72 net82 vgnd sky130_fd_io__refgen_res_ntwk_c
XR<4> net82 vcc_io_0p5 vgnd sky130_fd_io__refgen_res_ntwk_d
XR<5> vcc_io_0p5 net84 vgnd sky130_fd_io__refgen_res_ntwk_g
XR<6> net84 net153 vgnd sky130_fd_io__refgen_res_ntwk_h
XR<7> net153 net149 vgnd sky130_fd_io__refgen_res_ntwk_i
XI326 ibuf_sel_h_n in_lpf vinref vcc_a vgnd sky130_fd_io__refgen_in_lpf
XI343 ibuf_sel_h_n ibuf_sel_h net101 vcc_io vgnd sky130_fd_io__refgen_ls
XMP net76 net101 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=10 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRI340 net143 net146 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI339 net140 net143 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI338 net137 net140 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI337 net134 net137 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI336 vgnd net134 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI6 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=24.395
XRI335 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI334 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI333 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI332 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI331 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI330 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XRI11 vcc_io vcc_io vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=18.075
XI489 net153 sel_vcc_io_0p4 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI511 net149 sel_vcc_io vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_in_csw2 in out sel vcc_io vgnd
*.PININFO in:I sel:I vcc_io:I vgnd:I out:B
Xinv_vcc_io sel net24 vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x1
XI459 in net24 out vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI460 out sel in vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_in_csw in out sel vcc_io vgnd
*.PININFO in:I sel:I vcc_io:I vgnd:I out:B
Xinv_vcc_io sel net21 vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x1
XI460 out sel in vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI459 in net21 out vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI543 in sel vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_in_csw_vcc_io in out sel vcc_io vgnd
*.PININFO in:I sel:I vcc_io:I vgnd:I out:B
Xinv_vcc_io sel net35 vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x1
XI12 net49 out sky130_fd_io__refgen_em1o
XI66 in net27 sky130_fd_io__refgen_em1o
XI13 net27 vcc_io sky130_fd_io__refgen_em1s
XI14 net49 vcc_io sky130_fd_io__refgen_em1s
XI460 out sel in vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI459 net27 net35 net49 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI543 vcc_io vcc_io vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 vcc_io vcc_io net49 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_in_cswblk sel_vcc_io sel_vohref sel_vohref_0p5 vcc_io 
+ vcc_io_ref vgnd vinref_int vohref vohref_0p5 vohref_int
*.PININFO sel_vcc_io:I sel_vohref:I sel_vohref_0p5:I vcc_io_ref:I vgnd:I 
*.PININFO vohref:I vohref_0p5:I vohref_int:I vinref_int:O vcc_io:B
XI531 net51 net70 net53 vcc_io vgnd sky130_fd_io__refgen_in_csw2
XI517 net47 vinref_int sel_vohref vcc_io vgnd sky130_fd_io__refgen_in_csw
XI520 vohref_0p5 vinref_int sel_vohref_0p5 vcc_io vgnd sky130_fd_io__refgen_in_csw
XI514 vcc_io_ref vinref_int sel_vcc_io vcc_io vgnd 
+ sky130_fd_io__refgen_in_csw_vcc_io
XI9 net53 sel_vohref sky130_fd_io__refgen_em1o
XE1 net51 vohref sky130_fd_io__refgen_em1o
XE2 net70 vinref_int sky130_fd_io__refgen_em1s
XE0 net47 vohref_int sky130_fd_io__refgen_em1s
XI8 net53 vcc_io sky130_fd_io__refgen_em1s
.ENDS

.SUBCKT sky130_fd_io__refgen_in_xgates en_inpop_h fb_in fb_out ibuf_sel_h 
+ ibuf_sel_h_n ngate sel_vcc_io sel_vcc_io_0p4 sel_vohref sel_vohref_0p5 vcc_a 
+ vcc_io vgnd vinref vohref vohref_0p5
*.PININFO en_inpop_h:I fb_in:I ibuf_sel_h:I ibuf_sel_h_n:I ngate:I 
*.PININFO sel_vcc_io:I sel_vcc_io_0p4:I sel_vohref:I sel_vohref_0p5:I vohref:I 
*.PININFO vohref_0p5:I fb_out:O vinref:O vcc_a:B vcc_io:B vgnd:B
Xopamp en_inpop_h ibuf_sel_h_n fb_in vohref ngate fb_out vcc_a vgnd 
+ sky130_fd_io__refgen_opamp_stage_1
Xres_ntwk ibuf_sel_h ibuf_sel_h_n net57 sel_vcc_io sel_vcc_io_0p4 vcc_a vcc_io 
+ vcc_io_ref vgnd vinref sky130_fd_io__refgen_res_ntwk_vinref_1
Xcswblk sel_vcc_io sel_vohref sel_vohref_0p5 vcc_a vcc_io_ref vgnd net57 
+ vohref vohref_0p5 fb_out sky130_fd_io__refgen_in_cswblk
.ENDS

.SUBCKT sky130_fd_io__refgen_nor in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI3 net17 in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out in1 net17 vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 out in1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_inv_x2 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_in_logic en_inpop_h en_outop_h en_outop_h_n ibuf_sel_h 
+ ibuf_sel_h_n sel_vcc_io sel_vcc_io_0p4 sel_vohref sel_vohref_0p5 vcc_io vgnd 
+ vref_sel_h vref_sel_h_n vreg_en_h vtrip_sel_h vtrip_sel_h_n
*.PININFO ibuf_sel_h:I ibuf_sel_h_n:I vref_sel_h:I vref_sel_h_n:I vreg_en_h:I 
*.PININFO vtrip_sel_h:I vtrip_sel_h_n:I en_inpop_h:O en_outop_h:O 
*.PININFO en_outop_h_n:O sel_vcc_io:O sel_vcc_io_0p4:O sel_vohref:O 
*.PININFO sel_vohref_0p5:O vcc_io:B vgnd:B
XI488 vref_sel_h_n vtrip_sel_h net126 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI484 vref_sel_h vtrip_sel_h_n net119 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI483 net119 ibuf_sel_h sel_vohref_0p5 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI487 net126 ibuf_sel_h sel_vcc_io_0p4 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI485 vref_sel_h vtrip_sel_h net98 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI486 net98 ibuf_sel_h sel_vohref vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI482 vref_sel_h ibuf_sel_h sel_vcc_io vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nand2
XI439 vreg_en_h net70 net77 vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_nor
XI497 ibuf_sel_h_n vref_sel_h_n net70 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__refgen_nor
XI499 sel_vcc_io en_inpop_h vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x1
XI494 net77 en_outop_h vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x1
XI500 en_outop_h en_outop_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_inv_x2
.ENDS

.SUBCKT sky130_fd_io__refgen_in biasen_n en_outop_h en_outop_h_n fb_in fb_out 
+ hld_h_n hld_i_h_n hld_i_vpwr ibuf_sel ibuf_sel_h_n ngate od_h sel_vohref_0p5 
+ vcc_a vcc_io vgnd vinref vohref vohref_0p5 vpb vpwr vpwr_ka vref_sel vreg_en 
+ vtrip_sel
*.PININFO fb_in:I hld_h_n:I ibuf_sel:I ngate:I od_h:I vohref:I vohref_0p5:I 
*.PININFO vref_sel:I vreg_en:I vtrip_sel:I biasen_n:O en_outop_h:O 
*.PININFO en_outop_h_n:O fb_out:O hld_i_h_n:O hld_i_vpwr:O ibuf_sel_h_n:O 
*.PININFO sel_vohref_0p5:O vinref:O vcc_a:B vcc_io:B vgnd:B vpb:B vpwr:B 
*.PININFO vpwr_ka:B
Xxlators biasen_n hld_h_n hld_i_h_n hld_i_vpwr ibuf_sel ibuf_sel_h 
+ ibuf_sel_h_n en_outop_h en_outop_h_n od_h vcc_a vcc_io vgnd vpb vpwr vpwr_ka 
+ vref_sel vref_sel_h vref_sel_h_n vreg_en vreg_en_h net100 vtrip_sel 
+ vtrip_sel_h vtrip_sel_h_n sky130_fd_io__refgen_in_xlators
Xtransmission_gates en_inpop_h fb_in fb_out ibuf_sel_h ibuf_sel_h_n ngate 
+ sel_vcc_io sel_vcc_io_0p4 sel_vohref sel_vohref_0p5 vcc_a vcc_io vgnd vinref 
+ vohref vohref_0p5 sky130_fd_io__refgen_in_xgates
Xlogic en_inpop_h en_outop_h en_outop_h_n ibuf_sel_h ibuf_sel_h_n sel_vcc_io 
+ sel_vcc_io_0p4 sel_vohref sel_vohref_0p5 vcc_a vgnd vref_sel_h vref_sel_h_n 
+ vreg_en_h vtrip_sel_h vtrip_sel_h_n sky130_fd_io__refgen_in_logic
.ENDS

.SUBCKT sky130_fd_io__refgen_res_ntwk_a fb_out res_tap<8> res_tap<7> res_tap<6> 
+ res_tap<5> res_tap<4> res_tap<3> res_tap<2> res_tap<1> resgnd vgnd vohref_0p5
*.PININFO res_tap<8>:O res_tap<7>:O res_tap<6>:O res_tap<5>:O res_tap<4>:O 
*.PININFO res_tap<3>:O res_tap<2>:O res_tap<1>:O vohref_0p5:O fb_out:B 
*.PININFO resgnd:B vgnd:B
RI80 res_tap<8> fb_out sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
XRI0<17> int1<1> resgnd vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<16> int1<2> int1<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<15> int1<3> int1<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<14> int1<4> int1<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<13> int1<5> int1<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<12> int1<6> int1<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<11> int1<7> int1<6> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<10> int1<8> int1<7> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<9> int1<9> int1<8> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<8> int1<10> int1<9> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<7> int1<11> int1<10> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<6> int1<12> int1<11> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<5> int1<13> int1<12> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<4> int1<14> int1<13> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<3> int1<15> int1<14> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<2> int1<16> int1<15> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<1> int1<17> int1<16> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI0<0> res_tap<1> int1<17> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI68<1> int3 res_tap<21> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI68<0> res_tap<3> int3 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI63 res_tap<21> net63 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI62 res_tap<21> net63 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI61 res_tap<2> res_tap<11> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI60 res_tap<2> res_tap<11> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI59 res_tap<2> res_tap<11> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI58 res_tap<2> res_tap<11> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI65 net63 res_tap<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI66 net63 res_tap<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI64 net63 res_tap<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI67 net63 res_tap<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<8> int2<1> res_tap<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<7> int2<2> int2<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<6> int2<3> int2<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<5> int2<4> int2<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<4> int2<5> int2<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<3> int2<6> int2<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<2> int2<7> int2<6> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<1> int2<8> int2<7> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI50<0> res_tap<11> int2<8> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI69 net54 res_tap<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI71 vohref_0p5 net54 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI72 vohref_0p5 net54 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI73 res_tap<41> vohref_0p5 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI74 res_tap<41> vohref_0p5 vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<6> int5<1> res_tap<41> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<5> int5<2> int5<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<4> int5<3> int5<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<3> int5<4> int5<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<2> int5<5> int5<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<1> int5<6> int5<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI75<0> res_tap<5> int5<6> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI76<5> int4<1> res_tap<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI76<4> int4<2> int4<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI76<3> int4<3> int4<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI76<2> int4<4> int4<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI76<1> int4<5> int4<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI76<0> res_tap<4> int4<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI77<4> int6<1> res_tap<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI77<3> int6<2> int6<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI77<2> int6<3> int6<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI77<1> int6<4> int6<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI77<0> res_tap<6> int6<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<9> int7<1> res_tap<6> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<8> int7<2> int7<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<7> int7<3> int7<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<6> int7<4> int7<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<5> int7<5> int7<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<4> int7<6> int7<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<3> int7<7> int7<6> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<2> int7<8> int7<7> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<1> int7<9> int7<8> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI78<0> res_tap<7> int7<9> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<14> int8<1> res_tap<7> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<13> int8<2> int8<1> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<12> int8<3> int8<2> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<11> int8<4> int8<3> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<10> int8<5> int8<4> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<9> int8<6> int8<5> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<8> int8<7> int8<6> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<7> int8<8> int8<7> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<6> int8<9> int8<8> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<5> int8<10> int8<9> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<4> int8<11> int8<10> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<3> int8<12> int8<11> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<2> int8<13> int8<12> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<1> int8<14> int8<13> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
XRI79<0> res_tap<8> int8<14> vgnd sky130_fd_pr__res_generic_nd m=1 w=0.5 l=6.465
.ENDS

.SUBCKT sky130_fd_io__refgen_out_resblk fb_out res_stack res_tap<7> res_tap<6> 
+ res_tap<5> res_tap<4> res_tap<3> res_tap<2> res_tap<1> res_tap<0> 
+ sel_vohref_0p5 vcc vgnd vnb vohref_0p5
*.PININFO sel_vohref_0p5:I vcc:I vgnd:I vnb:I res_tap<7>:O res_tap<6>:O 
*.PININFO res_tap<5>:O res_tap<4>:O res_tap<3>:O res_tap<2>:O res_tap<1>:O 
*.PININFO res_tap<0>:O vohref_0p5:O fb_out:B res_stack:B
XI11 res_stack net40<0> net40<1> net40<2> net40<3> net40<4> net40<5> net40<6> 
+ net40<7> net041 vgnd vohref_0p5 sky130_fd_io__refgen_res_ntwk_a
XI10 fb_out res_tap<7> res_tap<6> res_tap<5> res_tap<4> res_tap<3> res_tap<2> 
+ res_tap<1> res_tap<0> vgnd vgnd net41 sky130_fd_io__refgen_res_ntwk_a
XI19 net041 sel_vohref_0p5 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=7 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_opamp_stage en_outop_h_n ibuf_sel_h_n inn inp ngate 
+ out vcc vcc_virt_i vcc_virt_o vgnd
*.PININFO en_outop_h_n:I ibuf_sel_h_n:I inn:I inp:I vcc:I vgnd:I out:O 
*.PININFO vcc_virt_i:O vcc_virt_o:O ngate:B
XI153 net140 vsource sky130_fd_io__refgen_em1o
XI220 net144 vsource sky130_fd_io__refgen_em1o
XI223 net136 vsource sky130_fd_io__refgen_em1o
XI214 net156 net97 sky130_fd_io__refgen_em1o
XI211 net156 net59 sky130_fd_io__refgen_em1o
XI215 vcc_virt_o net97 sky130_fd_io__refgen_em1s
XI212 vcc_virt_o net59 sky130_fd_io__refgen_em1s
XI227 vcc_virt_o en_outop_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI232 vcc_virt_i ibuf_sel_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI229 vcc_virt_o en_outop_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<1> out net59 vcc_virt_o vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI226 vcc_virt_o en_outop_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<2> net156 net156 vcc_virt_o vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<0> net156 net97 vcc_virt_o vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI228 vcc_virt_o en_outop_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP<3> out net156 vcc_virt_o vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI233 vcc_virt_i ibuf_sel_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI237 vcc_virt_i ibuf_sel_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI236 vcc_virt_i ibuf_sel_h_n vcc vcc sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI217<3> vcc_virt_o vcc_virt_o vcc_virt_o vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI216<3> vcc_virt_o vcc_virt_o vcc_virt_o vcc sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> vsource ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM<2> net144 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> net140 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM<3> net136 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI240<1> vsource vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI219 out vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN2 out inn vsource vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1 net156 inp vsource vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI218 net156 vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_opamp_biasgen_1 biasen_n ngate vgnd vpwr_ka
*.PININFO biasen_n:I vgnd:I vpwr_ka:I ngate:B
XI330 ngate net100 sky130_fd_io__refgen_em1o
XI235 net111 net113 sky130_fd_io__refgen_em1o
XI337 ngate net0166 sky130_fd_io__refgen_em1o
XI234 ngate net111 sky130_fd_io__refgen_em1o
XI187 net113 biasen_n vpwr_ka vpwr_ka sky130_fd_pr__pfet_01v8 m=2 w=5.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI334 ngate biasen_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> net100 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMopt net0166 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> ngate ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XRI298 net236 net111 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI299 net234 net236 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI300 net232 net234 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI301 net230 net232 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI302 net229 net230 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI303 net227 net228 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI304 net228 net226 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI305 net226 net224 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI306 net224 net222 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI307 net222 net229 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI308 net216 net227 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI309 net214 net216 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI310 net212 net214 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI311 net210 net212 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI312 net209 net210 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI313 net207 net208 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI314 net208 net206 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI315 net206 net204 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI316 net204 net202 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI317 net202 net209 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI318 net196 net207 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI319 net194 net196 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI320 net192 net194 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI321 net190 net192 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI322 net189 net190 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI323 ngate net188 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI324 net188 net186 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI325 net186 net184 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI326 net184 net182 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI327 net182 net189 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI267 net176 net113 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI266 net174 net176 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI265 net172 net174 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI264 net170 net172 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI263 net169 net170 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI262 net167 net168 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI261 net168 net166 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI260 net166 net164 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI259 net164 net162 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI258 net162 net169 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI257 net156 net167 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI256 net154 net156 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI255 net152 net154 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI254 net150 net152 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI253 net149 net150 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI252 net147 net148 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI251 net148 net146 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI250 net146 net144 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI249 net144 net142 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI248 net142 net149 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI247 net136 net147 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI246 net134 net136 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI245 net132 net134 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI244 net130 net132 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI243 net129 net130 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI242 net111 net128 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI241 net128 net126 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI240 net126 net124 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI239 net124 net122 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI238 net122 net129 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
XRI237 net113 net113 sky130_fd_pr__res_generic_po m=1 w=0.33 l=18.68
.ENDS

.SUBCKT sky130_fd_io__refgen_opamp_1 biasen_n en_outop_h_n ibuf_sel_h_n inn inp 
+ ngate out vcc vcc_virt_i vcc_virt_o vgnd vpwr_ka
*.PININFO biasen_n:I en_outop_h_n:I ibuf_sel_h_n:I inn:I inp:I vcc:I vgnd:I 
*.PININFO vpwr_ka:I ngate:O out:O vcc_virt_i:O vcc_virt_o:O
XI192 ngate en_outop_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xopamp_stage en_outop_h_n ibuf_sel_h_n inn inp ngate out vcc vcc_virt_i 
+ vcc_virt_o vgnd sky130_fd_io__refgen_opamp_stage
Xbias_stage biasen_n ngate vgnd vpwr_ka sky130_fd_io__refgen_opamp_biasgen_1
.ENDS

.SUBCKT sky130_fd_io__refgen_out_sub_rc in mid out vgnd
*.PININFO in:I vgnd:I mid:B out:B
XI484 net44 mid sky130_fd_io__refgen_em1s
XI2 net56 in sky130_fd_io__refgen_em1s
XI81 net60 in sky130_fd_io__refgen_em1s
XI8 net54 in sky130_fd_io__refgen_em1s
XI5 net52 in sky130_fd_io__refgen_em1s
XI10 net58 in sky130_fd_io__refgen_em1s
XI13 net50 in sky130_fd_io__refgen_em1s
XI16 net48 in sky130_fd_io__refgen_em1s
XI80 net97 out sky130_fd_io__refgen_em1s
XI95 net100 out sky130_fd_io__refgen_em1s
XI94 net103 out sky130_fd_io__refgen_em1s
XI93 net109 out sky130_fd_io__refgen_em1s
XI92 net106 out sky130_fd_io__refgen_em1s
XI109 net091 in sky130_fd_io__refgen_em1s
XI108 net093 in sky130_fd_io__refgen_em1s
XI103 net095 in sky130_fd_io__refgen_em1s
XI99 net097 in sky130_fd_io__refgen_em1s
XI82 net60 vgnd sky130_fd_io__refgen_em1o
XI9 net58 vgnd sky130_fd_io__refgen_em1o
XI1 net56 vgnd sky130_fd_io__refgen_em1o
XI7 net54 vgnd sky130_fd_io__refgen_em1o
XI6 net52 vgnd sky130_fd_io__refgen_em1o
XI14 net50 vgnd sky130_fd_io__refgen_em1o
XI15 net48 vgnd sky130_fd_io__refgen_em1o
XI73 net97 mid sky130_fd_io__refgen_em1o
XI72 net44 out sky130_fd_io__refgen_em1o
XI74 net109 mid sky130_fd_io__refgen_em1o
XI75 net100 mid sky130_fd_io__refgen_em1o
XI76 net94 out sky130_fd_io__refgen_em1o
XI111 net091 vgnd sky130_fd_io__refgen_em1o
XI110 net093 vgnd sky130_fd_io__refgen_em1o
XI104 net095 vgnd sky130_fd_io__refgen_em1o
XI100 net097 vgnd sky130_fd_io__refgen_em1o
XRI88 net106 net109 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=21.71
XRI79 net97 net106 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=21.71
XRI89 net109 net103 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=21.71
XRI90 net103 net100 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=21.71
XRI87 net94 net97 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=17.375
XRI24 net44 net94 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=17.375
XRI96 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=21.71
XRI91 out out vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.4 l=21.71
XI67 mid net60 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI483 mid net54 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 mid net56 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 mid net52 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 mid net58 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 mid net50 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 mid net48 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI117 mid net093 mid mid sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI113 mid net091 mid mid sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI112 mid net093 mid mid sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI105 mid net095 mid mid sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI116 mid net091 mid mid sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI115 mid net095 mid mid sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI101 mid net097 mid mid sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI114 mid net097 mid mid sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_out_sub en_outop_h en_outop_h_n fb_out pgate res_stack 
+ vcc_io vcc_virt_i vcc_virt_o vdda vgnd voutref
*.PININFO en_outop_h:I en_outop_h_n:I pgate:I vcc_io:I vcc_virt_i:I 
*.PININFO vcc_virt_o:I vdda:I vgnd:I fb_out:O res_stack:O voutref:O
Xrc_comp pgate mid voutref vgnd sky130_fd_io__refgen_out_sub_rc
XI70 pgate net94 sky130_fd_io__refgen_em1o
XI73 pgate net92 sky130_fd_io__refgen_em1o
XI42 net114 net90 sky130_fd_io__refgen_em1o
XI74 pgate net88 sky130_fd_io__refgen_em1o
XI9 net87 net133 sky130_fd_io__refgen_em1o
XI466 net85 net153 sky130_fd_io__refgen_em1o
XI43 net116 net82 sky130_fd_io__refgen_em1o
XI72 pgate net80 sky130_fd_io__refgen_em1o
XI87 voutref net193 sky130_fd_io__refgen_em1o
XI467 voutref net105 sky130_fd_io__refgen_em1s
XI40 net110 net116 sky130_fd_io__refgen_em1s
XI41 net112 net114 sky130_fd_io__refgen_em1s
XI39 net111 net112 sky130_fd_io__refgen_em1s
XI38 net111 net110 sky130_fd_io__refgen_em1s
XI28 voutref net103 sky130_fd_io__refgen_em1s
XI71 net80 vcc_io sky130_fd_io__refgen_em1s
XI29 net105 net85 sky130_fd_io__refgen_em1s
XI27 net103 net87 sky130_fd_io__refgen_em1s
XI75 net88 vcc_io sky130_fd_io__refgen_em1s
XI69 net94 vcc_io sky130_fd_io__refgen_em1s
XI76 net92 vcc_io sky130_fd_io__refgen_em1s
XI244 pgate en_outop_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> net105 pgate vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<7> net112 pgate vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<6> net110 pgate vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> net103 pgate vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<2> net85 pgate vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI13<5> vcc_virt_i vcc_virt_i vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=6 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI12<5> vcc_virt_o vcc_virt_o vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=6 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<11> net90 net88 vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<4> net153 net80 vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<9> net114 pgate vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<10> net82 net92 vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<8> net116 pgate vcc_virt_i vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<3> net87 pgate vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<5> net133 net94 vcc_virt_o vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=7.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1<5> voutref voutref fb_out fb_out sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1<4> voutref voutref fb_out fb_out sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1<3> voutref voutref fb_out fb_out sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1<2> voutref voutref fb_out fb_out sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1<1> voutref voutref fb_out fb_out sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1<0> voutref voutref fb_out fb_out sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI454<5> net111 net111 res_stack res_stack sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI454<4> net111 net111 res_stack res_stack sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI454<3> net111 net111 res_stack res_stack sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI454<2> net111 net111 res_stack res_stack sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI454<1> net111 net111 res_stack res_stack sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI454<0> net111 net111 res_stack res_stack sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI571 net193 en_outop_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_out biasen_n en_outop_h en_outop_h_n fb_in fb_out 
+ ibuf_sel_h_n ngate res_tap<7> res_tap<6> res_tap<5> res_tap<4> res_tap<3> 
+ res_tap<2> res_tap<1> res_tap<0> sel_vohref_0p5 vcc_io vdda vgnd vnb vohref 
+ vohref_0p5 voutref vpwr_ka
*.PININFO biasen_n:I en_outop_h:I en_outop_h_n:I fb_in:I ibuf_sel_h_n:I 
*.PININFO sel_vohref_0p5:I vohref:I fb_out:O ngate:O res_tap<7>:O res_tap<6>:O 
*.PININFO res_tap<5>:O res_tap<4>:O res_tap<3>:O res_tap<2>:O res_tap<1>:O 
*.PININFO res_tap<0>:O voutref:O vcc_io:B vdda:B vgnd:B vnb:B vohref_0p5:B 
*.PININFO vpwr_ka:B
Xresblk fb_out net41 res_tap<7> res_tap<6> res_tap<5> res_tap<4> res_tap<3> 
+ res_tap<2> res_tap<1> res_tap<0> sel_vohref_0p5 vcc_io vgnd vnb vohref_0p5 
+ sky130_fd_io__refgen_out_resblk
Xopamp biasen_n en_outop_h_n ibuf_sel_h_n vohref fb_in ngate net60 vcc_io 
+ net54 net55 vgnd vpwr_ka sky130_fd_io__refgen_opamp_1
Xrefgen_out_sub en_outop_h en_outop_h_n fb_out net60 net41 vcc_io net54 net55 
+ vdda vgnd voutref sky130_fd_io__refgen_out_sub
.ENDS

.SUBCKT sky130_fd_io__refgen_ref_mux amuxbus_a amuxbus_b sel_vdda_amuxbusa 
+ sel_vdda_amuxbusb sel_vdda_vref sel_vddio_amuxbusa sel_vddio_amuxbusb 
+ sel_vddio_vref vdda vohref vref vssa vswitch
*.PININFO amuxbus_a:I amuxbus_b:I sel_vdda_amuxbusa:I sel_vdda_amuxbusb:I 
*.PININFO sel_vdda_vref:I sel_vddio_amuxbusa:I sel_vddio_amuxbusb:I 
*.PININFO sel_vddio_vref:I vref:I vohref:O vdda:B vssa:B vswitch:B
XI39 vref vohref sel_vdda_vref sel_vddio_vref vdda vssa vswitch 
+ sky130_fd_io__refgen_t_switch
XI43 amuxbus_a vohref sel_vdda_amuxbusa sel_vddio_amuxbusa vdda vssa vswitch 
+ sky130_fd_io__refgen_t_switch
XI44 amuxbus_b vohref sel_vdda_amuxbusb sel_vddio_amuxbusb vdda vssa vswitch 
+ sky130_fd_io__refgen_t_switch
.ENDS

.SUBCKT sky130_fd_io__refgen_compl_switch in out sel vcc_io vgnd vnb
*.PININFO in:I sel:I out:O vcc_io:B vgnd:B vnb:B
XI114 sel sel_b vgnd vgnd vcc_io vcc_io sky130_fd_io__refgen_hvsbt_inv_x1
XI1 out sel_b in vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=5 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 in sel out vgnd sky130_fd_pr__nfet_g5v0d10v5 m=5 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__refgen_mux_top fb_in in<7> in<6> in<5> in<4> in<3> in<2> 
+ in<1> in<0> sel<7> sel<6> sel<5> sel<4> sel<3> sel<2> sel<1> sel<0> vddio 
+ vssio
*.PININFO in<7>:I in<6>:I in<5>:I in<4>:I in<3>:I in<2>:I in<1>:I in<0>:I 
*.PININFO sel<7>:I sel<6>:I sel<5>:I sel<4>:I sel<3>:I sel<2>:I sel<1>:I 
*.PININFO sel<0>:I fb_in:O vddio:B vssio:B
XI92 in<2> fb_in sel<5> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI90 in<4> fb_in sel<3> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI94 in<0> fb_in sel<7> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI9 in<7> fb_in sel<0> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI88 in<6> fb_in sel<1> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI89 in<5> fb_in sel<2> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI93 in<1> fb_in sel<6> vddio vssio vssio sky130_fd_io__refgen_compl_switch
XI91 in<3> fb_in sel<4> vddio vssio vssio sky130_fd_io__refgen_compl_switch
.ENDS

.SUBCKT sky130_fd_io__top_refgen_new amuxbus_a amuxbus_b dft_refgen enable_h 
+ enable_vdda_h hld_h_n ibuf_sel refleak_bias vccd vcchib vdda vddio vddio_q 
+ vinref vinref_dft voh_sel<2> voh_sel<1> voh_sel<0> vohref voutref 
+ voutref_dft vref_sel<1> vref_sel<0> vreg_en vssa vssd vssio vssio_q vswitch 
+ vtrip_sel
*.PININFO dft_refgen:I enable_h:I enable_vdda_h:I hld_h_n:I ibuf_sel:I 
*.PININFO voh_sel<2>:I voh_sel<1>:I voh_sel<0>:I vohref:I vref_sel<1>:I 
*.PININFO vref_sel<0>:I vreg_en:I vtrip_sel:I vinref:O voutref:O amuxbus_a:B 
*.PININFO amuxbus_b:B refleak_bias:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B 
*.PININFO vinref_dft:B voutref_dft:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
XI248 dft_refgen dft_refgen_vdda_n dft_refgen_vswitch enable_h enable_vdda_h 
+ hld_i_h_n hld_i_vpwr od_h sel_fb_mux<7> sel_fb_mux<6> sel_fb_mux<5> 
+ sel_fb_mux<4> sel_fb_mux<3> sel_fb_mux<2> sel_fb_mux<1> sel_fb_mux<0> 
+ net0106 net0105 net0104 net0103 net0102 net0101 vccd vdda vddio_q voh_sel<2> 
+ voh_sel<1> voh_sel<0> vref_sel<1> vref_sel<0> vref_sel_int vssa vssd vswitch 
+ sky130_fd_io__refgen_ctl
XI247 dft_refgen_vdda_n dft_refgen_vswitch vdda vinref vinref_dft voutref 
+ voutref_dft vssa vswitch sky130_fd_io__refgen_dft
Xrefgen_in biasen_n en_outop_h en_outop_h_n fb_vinref fb_vinref hld_h_n 
+ hld_i_h_n hld_i_vpwr ibuf_sel ibuf_sel_h_n refleak_bias od_h sel_vohref_0p5 
+ vddio_q vddio_q vssd vinref vohref_int vohref_0p5 vccd vccd vcchib 
+ vref_sel_int vreg_en vtrip_sel sky130_fd_io__refgen_in
Xrefgen_out biasen_n en_outop_h en_outop_h_n fb net88 ibuf_sel_h_n 
+ refleak_bias res_tap<7> res_tap<6> res_tap<5> res_tap<4> res_tap<3> 
+ res_tap<2> res_tap<1> res_tap<0> sel_vohref_0p5 vddio_q vdda vssd vssd 
+ vohref_int vohref_0p5 voutref vcchib sky130_fd_io__refgen_out
XI44 amuxbus_a amuxbus_b net0106 net0105 net0104 net0103 net0102 net0101 vdda 
+ vohref_int vohref vssa vswitch sky130_fd_io__refgen_ref_mux
XI43 fb res_tap<7> res_tap<6> res_tap<5> res_tap<4> res_tap<3> res_tap<2> 
+ res_tap<1> res_tap<0> sel_fb_mux<7> sel_fb_mux<6> sel_fb_mux<5> 
+ sel_fb_mux<4> sel_fb_mux<3> sel_fb_mux<2> sel_fb_mux<1> sel_fb_mux<0> 
+ vswitch vssa sky130_fd_io__refgen_mux_top
.ENDS

.SUBCKT sky130_fd_io__sio_gpio_in_buf en_h in_h in_vt out_h out_h_n vcc_io vgnd 
+ vpwr vtrip_sel_h_n
*.PININFO en_h:I in_h:I in_vt:I vcc_io:I vgnd:I vpwr:I vtrip_sel_h_n:I out_h:O 
*.PININFO out_h_n:O
Xttl_pd_op net82 net106 sky130_fd_io__tk_em1o
XI576 vtrip_sel_h_n vtrip_sel_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xpd2 net122 out_a vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1_mid_nat net118 vpwr net95 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpd_hrng net106 in_vt net105 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=3.00 l=1.00 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpden_1 net105 en_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpd1 net106 in_h net105 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI598 net106 out_a vcc_io vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI592 out_h out_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI584 net95 net95 out_a vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI571 net106 out_a vcc_io vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI597 net106 out_a net125 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI574 net106 out_a net125 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI570 out_a in_h net106 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI595 net82 in_vt net105 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=3.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI589 out_h_n net122 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xdis_trip_sel1 in_vt vtrip_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu2 net122 out_a vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1 net157 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpuen_2 out_a en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1_midopt net157 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI567 net118 in_h net157 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI568 vgnd out_a net157 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI590 out_h_n net122 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI579 net141 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI578 out_a in_h net141 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI593 out_h out_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI577 out_a vtrip_sel_h net118 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI582 vgnd out_a net141 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI575 vcc_io vtrip_sel_h net125 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_inbuf_ls en_h in_c in_t out_c out_t vgnd vpb vpwr
*.PININFO en_h:I in_c:I in_t:I vgnd:I vpb:I vpwr:I out_c:O out_t:O
XI534 out_t out_c vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_c out_t vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI536 out_c in_t vgnd_en vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_t in_c vgnd_en vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI552 vgnd_en en_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_inbuf_ls en en_h en_n in_c in_t out_ls vgnd vpb vpwr
*.PININFO en:I en_h:I en_n:I in_c:I in_t:I vgnd:I vpb:I vpwr:I out_ls:O
Xcom_ls en_h in_c in_t ls_out_n ls_out vgnd vpb vpwr 
+ sky130_fd_io__sio_com_inbuf_ls
XI561 ls_out_n en vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI54 ls_out en_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI44 ls_out_n out_ls vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 
+ psa=265e-3 pl=0.18 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=0.18 
+ nw=1.00 nm=1
.ENDS

.SUBCKT sky130_fd_io__sio_com_inbuf_einv ie ie_n in out vgnd vpb vpwr
*.PININFO ie:I ie_n:I in:I vgnd:I vpb:I vpwr:I out:O
XI2 out in n<1> vgnd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 n<1> ie vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in n<0> vpb sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 n<0> ie_n vpwr vpb sky130_fd_pr__pfet_01v8 m=2 w=5.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_inbuf_einv_hv ie ie_n in out vcc_io vgnd
*.PININFO ie:I ie_n:I in:I vcc_io:I vgnd:I out:O
XI2 out in n<1> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 n<1> ie vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in n<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 n<0> ie_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=6 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_inbuf_hvinv_x2 in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_inbuf_hvinv_x1 in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_inbuf en en_h en_h_n en_n ibufmux_out_h_n ibufmux_out_n 
+ in_h in_vt vcc_io vgnd vpb_ka vpwr_ka vtrip_sel_h_n
*.PININFO en:I en_h:I en_h_n:I en_n:I in_h:I in_vt:I vcc_io:I vgnd:I vpb_ka:I 
*.PININFO vpwr_ka:I vtrip_sel_h_n:I ibufmux_out_h_n:O ibufmux_out_n:O
Xbuf en_h in_h in_vt out_h_wo_buf out_h_n vcc_io vgnd vpwr_ka vtrip_sel_h_n 
+ sky130_fd_io__sio_gpio_in_buf
Xls en en_h en_n out_h_n out_h_wo_buf out_ls vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_inbuf_ls
Xen_lv_inv en en_n out_ls ibufmux_out_n vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_com_inbuf_einv
Xen_hv_inv en_h en_h_n out_h_buf ibufmux_out_h_n vcc_io vgnd 
+ sky130_fd_io__sio_com_inbuf_einv_hv
Xhv_inv_2x out_h_wo_buf_inv out_h_buf vcc_io vgnd vgnd 
+ sky130_fd_io__sio_inbuf_hvinv_x2
Xhv_inv_1x out_h_wo_buf out_h_wo_buf_inv vcc_io vgnd vgnd 
+ sky130_fd_io__sio_inbuf_hvinv_x1
.ENDS

.SUBCKT sky130_fd_io__sio_ibuf_se en en_h en_h_n en_n ibufmux_out_h_n ibufmux_out_n 
+ in_h in_vt vcc_io vgnd vpb_ka vpwr_ka vtrip_sel_h_n
*.PININFO en:I en_h:I en_h_n:I en_n:I in_h:I in_vt:I vcc_io:I vgnd:I vpb_ka:I 
*.PININFO vpwr_ka:I vtrip_sel_h_n:I ibufmux_out_h_n:O ibufmux_out_n:O
Xinbuf en en_h en_h_n en_n ibufmux_out_h_n ibufmux_out_n in_h in_vt vcc_io 
+ vgnd vpb_ka vpwr_ka vtrip_sel_h_n sky130_fd_io__sio_inbuf
.ENDS

.SUBCKT sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd gate in nbody nwellRing 
+ vgnd
*.PININFO gate:I in:B nbody:B nwellRing:B vgnd:B
XI1 in gate vgnd nbody sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=5.40 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.048 perim=0.94
RI9 net18 nbody sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI8 net16 nwellRing sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__sio_res250only_small_esd pad rout
*.PININFO pad:B rout:B
* XRI175 net12 net16 sky130_fd_pr__res_generic_po m=1 w=2 l=10.07
* XRI229 net16 rout sky130_fd_pr__res_generic_po m=1 w=2 l=0.17
* XRI228 pad net12 sky130_fd_pr__res_generic_po m=1 w=2 l=0.17
* RI237<1> net16 rout sky130_fd_pr__res_generic_m1
* RI237<2> net16 rout sky130_fd_pr__res_generic_li
* RI234<1> pad net12 sky130_fd_pr__res_generic_m1
* RI234<2> pad net12 sky130_fd_pr__res_generic_li

* NOTE: Removed all but the primary resistor;  the other devices do not
* show up in the layout.

XRI175 pad rout sky130_fd_pr__res_generic_po m=1 w=2 l=10.07
.ENDS

.SUBCKT sky130_fd_io__sio_buf_localesd in_h out_h out_vt vcc_io vgnd vtrip_sel_h
*.PININFO in_h:I vtrip_sel_h:I out_h:O out_vt:O vcc_io:B vgnd:B
Xggnfet2 vgnd out_vt vgnd vcc_io vgnd 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xggnfet6 vgnd vcc_io vgnd vcc_io out_h 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xggnfet5 vgnd vcc_io vgnd vcc_io out_vt 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xggnfet1 vgnd out_h vgnd vcc_io vgnd 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xesd_res in_h out_h sky130_fd_io__sio_res250only_small_esd
Xhv_passgate out_h vtrip_sel_h out_vt vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_inbuf_lv_dis ctl_in ctl_in_n din out vgnd vpb vpwr
*.PININFO ctl_in:I ctl_in_n:I din:I vgnd:I vpb:I vpwr:I out:O
XI549 out din vgnd vgnd sky130_fd_pr__nfet_01v8 m=5 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI558 n<0> ctl_in vpwr vpb sky130_fd_pr__pfet_01v8 m=4 w=5.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI550 out din n<0> vpb sky130_fd_pr__pfet_01v8 m=2 w=5.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI559 vpwr ctl_in_n din vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_inbuf_hv_dis ctl_in ctl_in_n din out vcc_io vgnd
*.PININFO ctl_in:I ctl_in_n:I din:I vcc_io:I vgnd:I out:O
XI549 out din vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI558 n<0> ctl_in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI550 out din n<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI559 vcc_io ctl_in_n din vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_ctl_ls_out in_c in_t out_c out_t vgnd vpb vpwr
*.PININFO in_c:I in_t:I vgnd:I vpb:I vpwr:I out_c:O out_t:O
XI35 out_c_n out_c vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 psa=265e-3 
+ pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 nw=1.00 nm=1
XI36 out_t_n out_t vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 psa=265e-3 
+ pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 nw=1.00 nm=1
XI536 out_t_n in_t vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_c_n in_c vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI534 out_c_n out_t_n vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_t_n out_c_n vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_ictl_outls_bank ie_diff_sel ie_diff_sel_h 
+ ie_diff_sel_h_n ie_diff_sel_n ie_se_sel ie_se_sel_h ie_se_sel_h_n 
+ ie_se_sel_n inp_dis_i inp_dis_i_h inp_dis_i_h_n inp_dis_i_n vgnd vpb_ka 
+ vpwr_ka
*.PININFO ie_diff_sel_h:I ie_diff_sel_h_n:I ie_se_sel_h:I ie_se_sel_h_n:I 
*.PININFO inp_dis_i_h:I inp_dis_i_h_n:I vgnd:I vpb_ka:I vpwr_ka:I 
*.PININFO ie_diff_sel:O ie_diff_sel_n:O ie_se_sel:O ie_se_sel_n:O inp_dis_i:O 
*.PININFO inp_dis_i_n:O
Xgpio_sel ie_se_sel_h_n ie_se_sel_h ie_se_sel_n ie_se_sel vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_in_ctl_ls_out
Xsio_sel ie_diff_sel_h_n ie_diff_sel_h ie_diff_sel_n ie_diff_sel vgnd vpb_ka 
+ vpwr_ka sky130_fd_io__sio_in_ctl_ls_out
Xbuf_dis inp_dis_i_h_n inp_dis_i_h inp_dis_i_n inp_dis_i vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_in_ctl_ls_out
.ENDS

.SUBCKT sky130_fd_io__sio_com_ictl_logic dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> 
+ dm_h_n<1> dm_h_n<0> ibuf_sel_h ibuf_sel_h_n ie_diff_sel_h ie_diff_sel_h_n 
+ ie_se_sel_h ie_se_sel_h_n inp_dis_h inp_dis_h_n inp_dis_i_h inp_dis_i_h_n 
+ tripsel_i_h tripsel_i_h_n vcc_io vgnd vtrip_sel_h
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO ibuf_sel_h:I ibuf_sel_h_n:I inp_dis_h:I inp_dis_h_n:I vcc_io:I 
*.PININFO vgnd:I vtrip_sel_h:I ie_diff_sel_h:O ie_diff_sel_h_n:O ie_se_sel_h:O 
*.PININFO ie_se_sel_h_n:O inp_dis_i_h:O inp_dis_i_h_n:O tripsel_i_h:O 
*.PININFO tripsel_i_h_n:O
XI18 inp_dis_i_h_n net107 net90 sky130_fd_io__tk_opti
XI8 inp_dis_i_h net102 net148 sky130_fd_io__tk_opti
Xinpdis_inv net148 net90 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
Xdm10nand_inv nand_dm01 and_dm01 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x1
Xibuf_diff_inv ie_diff_sel_h_n ie_diff_sel_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x1
Xibuf_se_inv ie_se_sel_h_n ie_se_sel_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x1
XI14 net120 net108 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI13 net71 net66 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI17 net107 net102 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
Xtripsel_inv tripsel_i_h_n tripsel_i_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x1
Xibuf_diff inp_dis_i_h_n ibuf_sel_h ie_diff_sel_h_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xibuf_se ibuf_sel_h_n inp_dis_i_h_n ie_se_sel_h_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xinpdis dm_buf_dis inp_dis_h_n net148 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xdm210 dm_h_n<2> and_dm01 dm_buf_dis vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xdm10 dm_h_n<1> dm_h_n<0> nand_dm01 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI11 dm_h<2> dm_h<1> net71 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI15 net66 net108 net107 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI12 dm_h<0> inp_dis_h net120 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xtripsel_nand ie_se_sel_h vtrip_sel_h tripsel_i_h_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
.ENDS

.SUBCKT sky130_fd_io__sio_ictl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> ibuf_sel_h ibuf_sel_h_n ie_diff_sel ie_diff_sel_h ie_diff_sel_h_n 
+ ie_diff_sel_n ie_se_sel ie_se_sel_h ie_se_sel_h_n ie_se_sel_n inp_dis_h 
+ inp_dis_h_n inp_dis_i inp_dis_i_h inp_dis_i_h_n inp_dis_i_n tripsel_i_h 
+ tripsel_i_h_n vcc_io vgnd vpb_ka vpwr_ka vtrip_sel_h
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO ibuf_sel_h:I ibuf_sel_h_n:I inp_dis_h:I inp_dis_h_n:I vcc_io:I 
*.PININFO vgnd:I vpb_ka:I vpwr_ka:I vtrip_sel_h:I ie_diff_sel:O 
*.PININFO ie_diff_sel_h:O ie_diff_sel_h_n:O ie_diff_sel_n:O ie_se_sel:O 
*.PININFO ie_se_sel_h:O ie_se_sel_h_n:O ie_se_sel_n:O inp_dis_i:O 
*.PININFO inp_dis_i_h:O inp_dis_i_h_n:O inp_dis_i_n:O tripsel_i_h:O 
*.PININFO tripsel_i_h_n:O
Xoutls_bank ie_diff_sel ie_diff_sel_h ie_diff_sel_h_n ie_diff_sel_n ie_se_sel 
+ ie_se_sel_h ie_se_sel_h_n ie_se_sel_n inp_dis_i inp_dis_i_h inp_dis_i_h_n 
+ inp_dis_i_n vgnd vpb_ka vpwr_ka sky130_fd_io__sio_com_ictl_outls_bank
Xlogic dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> ibuf_sel_h 
+ ibuf_sel_h_n ie_diff_sel_h ie_diff_sel_h_n ie_se_sel_h ie_se_sel_h_n 
+ inp_dis_h inp_dis_h_n inp_dis_i_h inp_dis_i_h_n tripsel_i_h tripsel_i_h_n 
+ vcc_io vgnd vtrip_sel_h sky130_fd_io__sio_com_ictl_logic
.ENDS

.SUBCKT sky130_fd_io__sio_ipath_com dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> ibuf_sel_h ibuf_sel_h_n ibufmux_out_h_n ibufmux_out_n ie_diff_sel 
+ ie_diff_sel_h ie_diff_sel_h_n ie_diff_sel_n inp_dis_h inp_dis_h_n out out_h 
+ pad vcc_io vgnd vpb_ka vpwr_ka vtrip_sel_h vtrip_sel_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO ibuf_sel_h:I ibuf_sel_h_n:I inp_dis_h:I inp_dis_h_n:I vcc_io:I 
*.PININFO vgnd:I vpb_ka:I vpwr_ka:I vtrip_sel_h:I vtrip_sel_h_n:I 
*.PININFO ie_diff_sel:O ie_diff_sel_h:O ie_diff_sel_h_n:O ie_diff_sel_n:O 
*.PININFO out:O out_h:O ibufmux_out_h_n:B ibufmux_out_n:B pad:B
Xibuf_se ie_se_sel ie_se_sel_h ie_se_sel_h_n ie_se_sel_n ibufmux_out_h_n 
+ ibufmux_out_n in_h in_vt vcc_io vgnd vpb_ka vpwr_ka tripsel_i_h_n 
+ sky130_fd_io__sio_ibuf_se
Xesd pad in_h in_vt vcc_io vgnd tripsel_i_h sky130_fd_io__sio_buf_localesd
Xmux_lv inp_dis_i inp_dis_i_n ibufmux_out_n out vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_com_inbuf_lv_dis
Xmux_hv inp_dis_i_h inp_dis_i_h_n ibufmux_out_h_n out_h vcc_io vgnd 
+ sky130_fd_io__sio_com_inbuf_hv_dis
Xcom_ictl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> ibuf_sel_h 
+ ibuf_sel_h_n ie_diff_sel ie_diff_sel_h ie_diff_sel_h_n ie_diff_sel_n 
+ ie_se_sel ie_se_sel_h ie_se_sel_h_n ie_se_sel_n inp_dis_h inp_dis_h_n 
+ inp_dis_i inp_dis_i_h inp_dis_i_h_n inp_dis_i_n tripsel_i_h tripsel_i_h_n 
+ vcc_io vgnd vpb_ka vpwr_ka vtrip_sel_h sky130_fd_io__sio_ictl
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_dlyblk in out1 out2 vgnd vpb_ka vpwr_ka
*.PININFO in:I vgnd:I vpb_ka:I vpwr_ka:I out1:O out2:O
Xe1 invout<2> out1 sky130_fd_io__sio_tk_em1o
XI43 invout<3> out1 sky130_fd_io__sio_tk_em1o
XI44 invout<4> out1 sky130_fd_io__sio_tk_em1o
XI45 invout<5> out1 sky130_fd_io__sio_tk_em1o
XI46 invout<6> out1 sky130_fd_io__sio_tk_em1o
XI49 invout<7> out1 sky130_fd_io__sio_tk_em1o
XI51 invout<6> out2 sky130_fd_io__sio_tk_em1o
XI52 invout<5> out2 sky130_fd_io__sio_tk_em1o
XI53 invout<4> out2 sky130_fd_io__sio_tk_em1o
XI54 invout<3> out2 sky130_fd_io__sio_tk_em1o
XI55 invout<2> out2 sky130_fd_io__sio_tk_em1o
XI56 invout<1> out2 sky130_fd_io__sio_tk_em1o
XI57 invout<1> in sky130_fd_io__sio_tk_em1o
XI42 invout<1> out1 sky130_fd_io__sio_tk_em1s
XI48 invout<7> out2 sky130_fd_io__sio_tk_em1s
XI58 int_sh2 invout<1> sky130_fd_io__sio_tk_em1s
XI59 int_sh1 invout<1> sky130_fd_io__sio_tk_em1s
XI8 int_sh2 in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI38 invout<7> invout<6> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI22 invout<2> invout<1> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI25 invout<3> invout<2> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 invout<4> invout<3> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 invout<6> invout<5> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 invout<5> invout<4> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI40 invout<7> invout<6> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 int_sh1 in vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI23 invout<2> invout<1> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 invout<6> invout<5> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 invout<5> invout<4> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI26 invout<4> invout<3> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 invout<3> invout<2> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_inbuf_einv ie ie_n in out vgnd vpb vpwr
*.PININFO ie:I ie_n:I in:I vgnd:I vpb:I vpwr:I out:O
XI2 out in n<1> vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 n<1> ie vgnd vgnd sky130_fd_pr__nfet_01v8 m=6 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in n<0> vpb sky130_fd_pr__pfet_01v8 m=3 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 n<0> ie_n vpwr vpb sky130_fd_pr__pfet_01v8 m=6 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_inbuf_einv_hv ie ie_n in out vcc_io vgnd
*.PININFO ie:I ie_n:I in:I vcc_io:I vgnd:I out:O
XI2 out in n<1> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 n<1> ie vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in n<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=2 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI9 n<0> ie_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=2 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__nor2_p in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
Xn0 out in0 vgnd vnb sky130_fd_pr__nfet_01v8 m=nm0 w=nw0 l=nl0 mult=1 sa=n0sa sb=n0sb sd=n0sd 
+ topography=normal area=0.063 perim=1.14
Xn1 out in1 vgnd vnb sky130_fd_pr__nfet_01v8 m=nm1 w=nw1 l=nl1 mult=1 sa=n1sa sb=n1sb sd=n1sd 
+ topography=normal area=0.063 perim=1.14
Xp1 out in1 int1 vpb sky130_fd_pr__pfet_01v8 m=pm1 w=pw1 l=pl1 mult=1 sa=p1sa sb=p1sb sd=p1sd 
+ topography=normal area=0.063 perim=1.14
Xp0 int1 in0 vpwr vpb sky130_fd_pr__pfet_01v8 m=pm0 w=pw0 l=pl0 mult=1 sa=p0sa sb=p0sb sd=p0sd 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_ctlblk ie_diff_dly_n ie_diff_n ie_diff_sel_h 
+ ie_diff_sel_h_n ie_diff_sel_n out_h_n out_hv out_lv out_n pcasc vcc_io vgnd 
+ vpb_ka vpwr_ka
*.PININFO ie_diff_sel_h:I ie_diff_sel_h_n:I ie_diff_sel_n:I out_hv:I out_lv:I 
*.PININFO pcasc:I vcc_io:I vgnd:I vpb_ka:I vpwr_ka:I ie_diff_dly_n:O 
*.PININFO ie_diff_n:O out_h_n:O out_n:O
XI33 int<8> int<7> ie_diff_dly_n vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_in_diff_dlyblk
Xen_lv_inv int<10> int<11> out_lv out_n vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_inbuf_einv
Xen_hv_inv ie_diff_sel_h ie_diff_sel_h_n out_hv out_h_n vcc_io vgnd 
+ sky130_fd_io__sio_inbuf_einv_hv
XI31 ie_diff_n int<6> sky130_fd_io__sio_tk_em1o
XI32 int<8> int<6> sky130_fd_io__sio_tk_em1o
XI48 vgnd int<2> sky130_fd_io__sio_tk_em1o
XI28 ie_diff_n int<7> sky130_fd_io__sio_tk_em1s
XI29 int<8> int<9> sky130_fd_io__sio_tk_em1s
XI19 ie_diff_sel_n ie_diff_dly_n int<10> vgnd vgnd vpb_ka vpwr_ka sky130_fd_io__nor2_p 
+ p0sd=280e-3 p0sb=795e-3 p0sa=795e-3 pl0=0.25 pw0=1.00 pm0=1 p1sd=280e-3 
+ p1sb=265e-3 p1sa=1.325 pl1=0.25 pw1=1.00 pm1=1 n1sd=280e-3 n1sb=265e-3 
+ n1sa=1.325 nl1=0.25 nw1=1.00 nm1=1 n0sd=280e-3 n0sb=795e-3 n0sa=795e-3 
+ nl0=0.25 nw0=1.00 nm0=1
XI35 int<10> int<11> vgnd vgnd vpb_ka vpwr_ka sky130_fd_io__inv_p psd=280e-3 psb=265e-3 
+ psa=795e-3 pl=0.25 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=795e-3 nl=0.25 
+ nw=1.00 nm=1
Xdiffseln_nfet int<1> ie_diff_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 
+ sa=20 sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 int<1> int<3> int<2> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 int<4> int<1> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=20 sb=20 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI9 int<5> int<4> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=20 sb=20 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI46 int<3> int<1> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.80 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 int<9> int<4> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.80 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 int<6> int<5> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.80 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI44 int<2> int<3> vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xdiffselhn_p int<0> ie_diff_sel_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 
+ sa=20 sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpcasc_p int<1> pcasc int<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 int<4> int<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI10 int<5> int<4> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI16 int<6> int<9> vpwr_ka vpb_ka sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xlvp1 int<9> int<6> vpwr_ka vpb_ka sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI47 int<3> int<1> vpwr_ka vpb_ka sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.80 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_res_3k r0 r1 vnb
*.PININFO vnb:I r0:B r1:B
XI241 r0 net14 sky130_fd_io__sio_tk_em1s
XI240 net22 r1 sky130_fd_io__sio_tk_em1o
XRI248 r0 net14 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.68 l=1.53
XRI238 net22 r1 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.68 l=1.53
XRI237 net14 net22 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.68 l=8.405
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_res_9k r0 r1 vnb
*.PININFO vnb:I r0:B r1:B
Xe4 net15 net13 sky130_fd_io__sio_tk_em1s
Xe2 net033 r1 sky130_fd_io__sio_tk_em1s
Xe1 net37 net19 sky130_fd_io__sio_tk_em1s
Xe3 net19 net15 sky130_fd_io__sio_tk_em1s
Xe7 net9 net033 sky130_fd_io__sio_tk_em1s
Xe6 net11 net9 sky130_fd_io__sio_tk_em1s
Xe5 net13 net11 sky130_fd_io__sio_tk_em1s
Xe8 r0 net37 sky130_fd_io__sio_tk_em1o
XRr8 net9 net033 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3
XRr7 net11 net9 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3
XRr6 net13 net11 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3
XRr4 net19 net15 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3
XRr3 net033 r1 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4
XRr5 net15 net13 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3
XRrbase r0 net37 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20
XRr2 net37 net19 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_res_40k r0 r1 vnb
*.PININFO vnb:I r0:B r1:B
Xe5 net56 net54 sky130_fd_io__sio_tk_em1o
Xe4 net38 net56 sky130_fd_io__sio_tk_em1o
Xe3 net60 net58 sky130_fd_io__sio_tk_em1o
Xe2 net62 net60 sky130_fd_io__sio_tk_em1o
Xe1 r0 net62 sky130_fd_io__sio_tk_em1o
Xe6 net54 net52 sky130_fd_io__sio_tk_em1o
Xe7 net34 net50 sky130_fd_io__sio_tk_em1o
Xe12 net50 net48 sky130_fd_io__sio_tk_em1o
Xe13 net48 net46 sky130_fd_io__sio_tk_em1o
Xe14 net32 net44 sky130_fd_io__sio_tk_em1o
Xe15 net44 net42 sky130_fd_io__sio_tk_em1o
Xe16 net42 r1 sky130_fd_io__sio_tk_em1o
Xe9 net52 net36 sky130_fd_io__sio_tk_em1s
Xe11 net46 net32 sky130_fd_io__sio_tk_em1s
Xe10 net36 net34 sky130_fd_io__sio_tk_em1s
Xe8 net58 net38 sky130_fd_io__sio_tk_em1s
Xe20 net053 vnb sky130_fd_io__sio_tk_em1s
Xe19 net051 vnb sky130_fd_io__sio_tk_em1s
Xe17 r0 net050 sky130_fd_io__sio_tk_em1s
XRdummy1 net050 net0140 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20.8
XRdummy2 net051 net053 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20.8
XRr15 net42 r1 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20.8
XRr14 net44 net42 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20.8
XRr13 net32 net44 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=7
XRr12 net46 net32 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=12.4
XRr11 net48 net46 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=10.4
XRr10 net50 net48 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8
XRr9 net34 net50 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=7
XRr8 net36 net34 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.4
XRr7 net52 net36 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8.4
XRr6 net54 net52 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=7
XRr5 net56 net54 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=8
XRr4 net38 net56 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=10.4
XRr3 net58 net38 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=12.4
XRr2 net60 net58 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=7
XRr16 net62 net60 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20.8
XRrbase r0 net62 vnb sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=20.8
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_sub ie_diff_n ie_diff_sel_h nbias out_a out_a_hv 
+ out_b out_b_hv pad_esd pcasc vcc_io vcc_ioq vgnd vinref
*.PININFO ie_diff_n:I ie_diff_sel_h:I out_a_hv:I out_b_hv:I vcc_io:I vcc_ioq:I 
*.PININFO vgnd:I vinref:I out_a:O out_b:O pcasc:O nbias:B pad_esd:B
XI1819 n1bb1r ndiffcom vgnd sky130_fd_io__sio_in_diff_res_3k
XI1818 n1aa1r ndiffcom vgnd sky130_fd_io__sio_in_diff_res_3k
Xe2 net112 ndiffcom sky130_fd_io__tk_em1s
XI1700 net125 out_a sky130_fd_io__tk_em1o
XI1693 net123 net238 sky130_fd_io__tk_em1o
XI1696 net121 out_b sky130_fd_io__tk_em1o
XI1706 net119 net243 sky130_fd_io__tk_em1o
XI1811 net117 vgnd sky130_fd_io__tk_em1o
Xe3 net262 net112 sky130_fd_io__tk_em1o
Xe1 net274 net112 sky130_fd_io__tk_em1o
XI1810 net111 vgnd sky130_fd_io__tk_em1o
Xr1b vcc_ioq n1aa vgnd sky130_fd_io__sio_in_diff_res_9k
XI1787 vcc_ioq n1bb vgnd sky130_fd_io__sio_in_diff_res_9k
Xrcasc vcc_ioq net134 vgnd sky130_fd_io__sio_in_diff_res_40k
XRI1725 vgnd vgnd sky130_fd_pr__res_generic_po m=1 w=0.33 l=5.685
Xpdummy2 n1bb vcc_ioq pcasc vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1690 net123 pcasc n1aa vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdummy3 n1bb vcc_ioq vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1709 net119 pcasc n1bb vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdummy1 n1aa vcc_ioq vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=2 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1704 net125 pcasc n1aa vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1699 net121 pcasc n1bb vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpcap2 vcc_ioq pcasc vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpcdis pcasc ie_diff_sel_h vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpcap1 vcc_ioq pcasc vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=10 w=3.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpl2a net238 pcasc n1aa vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpl2b out_b pcasc n1bb vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpl3b net243 pcasc n1bb vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.5 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpl3a out_a pcasc n1aa vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.5 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpbias1 net134 pcasc pcasc vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1776 n1bb out_b_hv n1bb2s vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1774 n1aa out_a_hv n1aa1s vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1777 n1aa out_b_hv n1aa2s vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1775 n1bb out_a_hv n1bb1s vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1808 vgnd vgnd net111 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffbias net112 nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=16 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1809 vgnd vgnd net117 vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
Xncap vgnd nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=4.00 mult=5 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1735 n1aa2s pad_esd ndiffcom vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 
+ sa=1.445 sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
Xn3bdis net243 ie_diff_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1736 n1bb1s vinref ndiffcom vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
Xcmlpa out_a out_a vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.80 mult=1 sa=1.345 sb=2.425 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xn2adis net238 ie_diff_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffref n1bb2s vinref n1bb1r vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 
+ sa=1.445 sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
Xndb1 net274 nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffin n1aa1s pad_esd n1aa1r vgnd sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 
+ sa=1.445 sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
Xclmpb out_b out_b vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.80 mult=1 sa=1.345 sb=2.425 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xndb2 net262 nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffref3 net243 net243 vgnd vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.50 mult=1 sa=1.045 
+ sb=2.605 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1823 vgnd nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1822 vgnd nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=16 w=3.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xn2bdis out_b ie_diff_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xn3adis out_a ie_diff_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffin3 out_a net243 vgnd vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.50 mult=1 sa=2.605 
+ sb=1.045 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1821 nbias nbias nbias vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffin2 net238 net238 vgnd vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.50 mult=1 sa=1.045 
+ sb=2.605 sd=280e-3 topography=normal area=0.063 perim=1.14
Xndiffref2 out_b net238 vgnd vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.50 mult=1 sa=2.605 
+ sb=1.045 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnbias1a pcasc nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1820 nbias nbias nbias vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_biasgen_res ie_diff_sel_n ngate vgnd vpwr
*.PININFO ie_diff_sel_n:I vgnd:I vpwr:I ngate:B
Xo4 net100 net108 sky130_fd_io__sio_tk_em1s
Xo2 net102 net106 sky130_fd_io__sio_tk_em1s
Xo1 net106 net104 sky130_fd_io__sio_tk_em1s
Xo3 net108 net102 sky130_fd_io__sio_tk_em1s
Xo5 net101 net100 sky130_fd_io__sio_tk_em1s
Xo6 net96 net101 sky130_fd_io__sio_tk_em1s
Xo7 net94 net96 sky130_fd_io__sio_tk_em1s
Xo8 net116 net94 sky130_fd_io__sio_tk_em1s
Xos2 net90 net92 sky130_fd_io__sio_tk_em1s
Xos1 net104 net90 sky130_fd_io__sio_tk_em1s
Xo23 ngate net88 sky130_fd_io__sio_tk_em1s
Xo21 net112 net121 sky130_fd_io__sio_tk_em1o
Xo13 net134 net136 sky130_fd_io__sio_tk_em1o
Xo12 net114 net134 sky130_fd_io__sio_tk_em1o
Xo15 net122 net132 sky130_fd_io__sio_tk_em1o
Xo18 net124 net130 sky130_fd_io__sio_tk_em1o
Xo17 net130 net128 sky130_fd_io__sio_tk_em1o
Xo16 net128 net132 sky130_fd_io__sio_tk_em1o
Xo19 net120 net124 sky130_fd_io__sio_tk_em1o
Xo14 net136 net122 sky130_fd_io__sio_tk_em1o
Xo20 net121 net120 sky130_fd_io__sio_tk_em1o
Xo10 net119 net118 sky130_fd_io__sio_tk_em1o
Xo9 net118 net116 sky130_fd_io__sio_tk_em1o
Xo11 net119 net114 sky130_fd_io__sio_tk_em1o
Xo22 net88 net112 sky130_fd_io__sio_tk_em1o
Xos3 net92 net110 sky130_fd_io__sio_tk_em1o
XRres10k8 net124 net130 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k10 net121 net120 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres2k9 net118 net116 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres2k8 net116 net94 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres2k4 net100 net108 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres2k3 net108 net102 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres10k5 net122 net132 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres2k6 net96 net101 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=6.43
XRres2k5 net101 net100 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres2k2 net102 net106 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres10k6 net128 net132 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k2 net134 net114 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k11 net112 net121 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k7 net130 net128 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres2k7 net94 net96 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=6.43
XRres2k10 net119 net118 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres10k3 net134 net136 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k1 net114 net119 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres2k1 net106 net104 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5.785
XRres10k4 net136 net122 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k9 net120 net124 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRdummy2 vpwr vpwr vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRdummy1 vpwr vpwr vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XReres1 net104 net90 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4
XRdummy3 vpwr vpwr vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XReres3 net92 net110 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=3.705
XRres10k13 ngate net88 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRres10k12 net88 net112 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XRdummy4 vgnd vgnd vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=25.315
XReres2 net90 net92 vgnd sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4
XI187 net110 ie_diff_sel_n vpwr vpwr sky130_fd_pr__pfet_01v8 m=2 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_biasgen ie_diff_sel_h_n ie_diff_sel_n ngate vcc_io vgnd 
+ vpwr
*.PININFO ie_diff_sel_h_n:I ie_diff_sel_n:I vcc_io:I vgnd:I vpwr:I ngate:B
XI235 ie_diff_sel_n nbias vgnd vpwr sky130_fd_io__sio_biasgen_res
XRI322 net_152 pbias vgnd sky130_fd_pr__res_generic_nd m=1 w=0.33 l=43.375
XRI300 vgnd fb vgnd sky130_fd_pr__res_generic_nd m=1 w=0.33 l=173.5
XI344 vpwr_3 vpwr_3 vpwr_2 vpwr_2 sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI345 vpwr_2 vpwr_2 vpwr_1 vpwr_1 sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 fb net_152 fb fb sky130_fd_pr__nfet_05v0_nvt m=8 w=10.0 l=0.90 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI326 ngate ie_diff_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XIdiff_p net_108 fb com vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI296 ngate ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI276 nbias nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI277 nbias ie_diff_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XIbiasn com nbias vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XIdiff_n pbias vpwr_1 com vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI343 vpwr_4 vpwr_4 vpwr_3 vpwr_3 sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI365 vgnd ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI356 pbias pbias pbias vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI355 net_108 net_108 net_108 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI346 vpwr_1 vpwr_1 vgnd vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI316 net1 ie_diff_sel_n vpwr vpwr sky130_fd_pr__pfet_01v8_lvt m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI285 fb pbias net1 vpwr sky130_fd_pr__pfet_01v8_lvt m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XIloadp1 net_108 net_108 net1 vpwr sky130_fd_pr__pfet_01v8_lvt m=4 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XIloadp2 pbias net_108 net1 vpwr sky130_fd_pr__pfet_01v8_lvt m=4 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI295 net_178 pbias net1 vpwr sky130_fd_pr__pfet_01v8_lvt m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI359 vpwr vpwr net_178 vpwr sky130_fd_pr__pfet_01v8_lvt m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI357 vpwr vpwr net1 vpwr sky130_fd_pr__pfet_01v8_lvt m=2 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI354 ngate ie_diff_sel_n net_178 net_178 sky130_fd_pr__pfet_01v8_lvt m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI358 vpwr vpwr fb vpwr sky130_fd_pr__pfet_01v8_lvt m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI347 vpwr_4 ie_diff_sel_n vpwr vpwr sky130_fd_pr__pfet_01v8 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_lsblk ie_diff_dly_n ie_diff_n ie_diff_sel_h 
+ ie_diff_sel_h_n in_a in_b out out_h vcc_io vgnd vpb vpwr
*.PININFO ie_diff_dly_n:I ie_diff_n:I ie_diff_sel_h:I ie_diff_sel_h_n:I in_a:I 
*.PININFO in_b:I vcc_io:I vgnd:I vpb:I vpwr:I out:O out_h:O
XI1661 hvout_n hvout vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1640 hvout hvout_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1642 hlsin outb net101 vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xlvp2 outb out vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xlvp1 out outb vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI427 out_h net134 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI741 net134 hvout vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1643 hlsinb hlsin vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1651 net101 ie_diff_dly_n vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=3 w=1.00 l=0.18 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1659 net122 hlsin vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1663 hvout hvout_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1662 hvout_n hvout vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1656 hvout ie_diff_sel_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1646 net106 hlsinb vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1473 out ie_diff_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xlvn1 out in_a vgnd vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1658 hvout_n ie_diff_sel_h net142 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1657 hvout ie_diff_sel_h net150 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1649 hlsinb hlsin vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1645 net150 vpwr net106 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xlvn2 outb in_b vgnd vgnd sky130_fd_pr__nfet_01v8 m=3 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1660 net142 vpwr net122 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1648 hlsin outb vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI742 net134 hvout vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI428 out_h net134 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1654 hlsin ie_diff_dly_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_localesd ng_ctl pad pad_sw0 vcc_io vcc_ioq vgnd
*.PININFO ng_ctl:I vcc_io:I vcc_ioq:I vgnd:I pad:B pad_sw0:B
XI1718 pad_sw0 net56 sky130_fd_io__sio_tk_em1s
Xpad_esd_res pad net56 sky130_fd_io__sio_res250only_small_esd
Xesdfet2 vgnd net56 vgnd vcc_io vgnd 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xesdfet1 vgnd vcc_ioq vgnd vcc_io net56 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xesdfet4 vgnd pad_sw0 vgnd vcc_io vgnd 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
Xesdfet3 vgnd vcc_ioq vgnd vcc_io pad_sw0 
+ sky130_fd_io__sio_signal_5_sym_hv_local_5term_esd
XI1727 net56 ng_ctl pad_sw0 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff_iclmp ie_diff_sel_h ie_diff_sel_h_n nbias ng_ctl 
+ vcc_ioq vgnd vinref
*.PININFO ie_diff_sel_h:I ie_diff_sel_h_n:I vcc_ioq:I vgnd:I vinref:I ng_ctl:O 
*.PININFO nbias:B
XI1821 net221 ng_ctl sky130_fd_io__sio_tk_em1o
XI1810 net121 net137 sky130_fd_io__sio_tk_em1o
XI1806 net77 net118 sky130_fd_io__sio_tk_em1o
XI1802 net95 vcc_ioq sky130_fd_io__sio_tk_em1o
XI1800 vgnd net93 sky130_fd_io__sio_tk_em1o
XI1795 net113 net79 sky130_fd_io__sio_tk_em1o
XI1789 pbias_nsw net110 sky130_fd_io__sio_tk_em1o
XI1815 net89 net108 sky130_fd_io__sio_tk_em1o
XI1814 net107 net177 sky130_fd_io__sio_tk_em1o
XI1787 pbias_nsw net104 sky130_fd_io__sio_tk_em1o
XI1784 pbias_nsw net146 sky130_fd_io__sio_tk_em1o
XI1822 ng_ctl net100 sky130_fd_io__sio_tk_em1s
XI1808 net139 net121 sky130_fd_io__sio_tk_em1s
XI1809 net139 net136 sky130_fd_io__sio_tk_em1s
XI1801 net95 ie_diff_sel_h_n sky130_fd_io__sio_tk_em1s
XI1799 net93 ie_diff_sel_h sky130_fd_io__sio_tk_em1s
XI1788 net110 vcc_ioq sky130_fd_io__sio_tk_em1s
XI1813 net89 net177 sky130_fd_io__sio_tk_em1s
XI1812 ng_ctl net107 sky130_fd_io__sio_tk_em1s
XI1786 net104 vcc_ioq sky130_fd_io__sio_tk_em1s
XI1811 ng_ctl net176 sky130_fd_io__sio_tk_em1s
XI1796 net113 vgnd sky130_fd_io__sio_tk_em1s
XI1797 net79 nbias sky130_fd_io__sio_tk_em1s
XI1805 net77 net137 sky130_fd_io__sio_tk_em1s
XI1783 net146 vcc_ioq sky130_fd_io__sio_tk_em1s
Xpcdis pbias_nsw net93 vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1741 vcc_ioq pbias_nsw pbias_nsw vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1817 net177 vinref net176 ng_ctl sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1732 net137 vinref net121 net139 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1793 net118 vinref net121 net139 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1792 vcc_ioq pbias_nsw vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1728 net190 pbias_nsw vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1790 net202 net110 vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1816 net108 vinref net107 ng_ctl sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1791 net197 net95 vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1782 vcc_ioq net146 pbias_nsw vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1785 net190 net104 vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1803 net137 vinref net136 net139 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1818 net177 vinref net107 ng_ctl sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1776 net202 pbias_nsw vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 
+ sb=20 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1820 net100 net93 vcc_ioq vcc_ioq sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1819 net221 net95 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1742 pbias_nsw net79 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1733 net77 net93 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1794 pbias_nsw net113 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1779 net206 net206 ng_ctl vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1780 net202 net202 ng_ctl vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1778 net197 net190 net206 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1781 net89 net93 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=20 sb=20 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1763 net190 net190 net139 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=1.445 
+ sb=2.625 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_diff ie_diff_dly_n ie_diff_n ie_diff_sel_h 
+ ie_diff_sel_h_n ie_diff_sel_n out out_h pad_esd pcasc vcc_io vcc_ioq vgnd 
+ vinref vpb vpwr
*.PININFO ie_diff_dly_n:I ie_diff_n:I ie_diff_sel_h:I ie_diff_sel_h_n:I 
*.PININFO ie_diff_sel_n:I vcc_io:I vcc_ioq:I vgnd:I vinref:I vpb:I vpwr:I 
*.PININFO out:O out_h:O pcasc:O pad_esd:B
Xsub ie_diff_n ie_diff_sel_h net104 n3a out_a_hv n2b out_b_hv pad_esd1 pcasc 
+ vcc_io vcc_ioq vgnd vinref sky130_fd_io__sio_in_diff_sub
XI1655 out_b_hv out_a_hv vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x4
XI1654 net71 out_b_hv vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI1656 out_h net71 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
Xbias ie_diff_sel_h_n ie_diff_sel_n net104 vcc_io vgnd vpwr 
+ sky130_fd_io__sio_biasgen
Xlsblk ie_diff_dly_n ie_diff_n ie_diff_sel_h ie_diff_sel_h_n n3a n2b out out_h 
+ vcc_ioq vgnd vpb vpwr sky130_fd_io__sio_in_diff_lsblk
XI1638 net95 pad_esd pad_esd1 vcc_io vcc_ioq vgnd 
+ sky130_fd_io__sio_in_diff_localesd
XI1640 ie_diff_sel_h ie_diff_sel_h_n net104 net95 vcc_ioq vgnd vinref 
+ sky130_fd_io__sio_in_diff_iclmp
.ENDS

.SUBCKT sky130_fd_io__sio_ibuf_diff_tsg4 ie_diff_sel_h ie_diff_sel_h_n 
+ ie_diff_sel_n out_h_n out_n pad_esd sio_diff_hyst_en_h vcc_io vcc_ioq vgnd 
+ vinref vpb_ka vpwr_ka
*.PININFO ie_diff_sel_h:I ie_diff_sel_h_n:I ie_diff_sel_n:I 
*.PININFO sio_diff_hyst_en_h:I vcc_io:I vcc_ioq:I vgnd:I vinref:I vpb_ka:I 
*.PININFO vpwr_ka:I out_h_n:O out_n:O pad_esd:B
Xctlblk ie_diff_dly_n ie_diff_n ie_diff_sel_h ie_diff_sel_h_n ie_diff_sel_n 
+ out_h_n out_hv out_lv out_n pcasc vcc_ioq vgnd vpb_ka vpwr_ka 
+ sky130_fd_io__sio_in_diff_ctlblk
Xdiff ie_diff_dly_n ie_diff_n ie_diff_sel_h ie_diff_sel_h_n ie_diff_sel_n 
+ out_lv out_hv pad_esd pcasc vcc_io vcc_ioq vgnd vinref vpb_ka vpwr_ka 
+ sky130_fd_io__sio_in_diff
.ENDS

.SUBCKT sky130_fd_io__sio_ipath_tsg4 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> ibuf_sel_h ibuf_sel_h_n inp_dis_h inp_dis_h_n out out_h pad 
+ sio_diff_hyst_en_h vcc_io vcc_ioq vgnd vinref vpb_ka vpwr_ka vtrip_sel_h 
+ vtrip_sel_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO ibuf_sel_h:I ibuf_sel_h_n:I inp_dis_h:I inp_dis_h_n:I 
*.PININFO sio_diff_hyst_en_h:I vcc_io:I vcc_ioq:I vgnd:I vinref:I vpb_ka:I 
*.PININFO vpwr_ka:I vtrip_sel_h:I vtrip_sel_h_n:I out:O out_h:O pad:B
Xcom_ipath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> ibuf_sel_h 
+ ibuf_sel_h_n out_h_n_einv out_n_einv ie_diff_sel ie_diff_sel_h 
+ ie_diff_sel_h_n ie_diff_sel_n inp_dis_h inp_dis_h_n out out_h pad vcc_ioq 
+ vgnd vpb_ka vpwr_ka vtrip_sel_h vtrip_sel_h_n sky130_fd_io__sio_ipath_com
Xsio_ibuf ie_diff_sel_h ie_diff_sel_h_n ie_diff_sel_n out_h_n_einv out_n_einv 
+ pad sio_diff_hyst_en_h vcc_io vcc_ioq vgnd vinref vpb_ka vpwr_ka 
+ sky130_fd_io__sio_ibuf_diff_tsg4
.ENDS

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x8 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=8 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XI1 out in vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=8 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_lvlp_inv_x4 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI1 out in vpwr vpb sky130_fd_pr__pfet_01v8_hvt m=4 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 out in vgnd vnb sky130_fd_pr__nfet_01v8 m=4 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_ctl_ls_out in_c in_t out_c out_t vgnd vpwr
*.PININFO in_c:I in_t:I vgnd:I vpwr:I out_c:O out_t:O
XI35 out_c_n out_c vgnd vgnd vpwr vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 
+ psa=265e-3 pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 
+ nw=1.00 nm=1
XI36 out_t_n out_t vgnd vgnd vpwr vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 
+ psa=265e-3 pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 
+ nw=1.00 nm=1
XI536 out_t_n in_t vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_c_n in_c vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI534 out_c_n out_t_n vpwr vpwr sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_t_n out_c_n vpwr vpwr sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_ctl_ls hld_h_n in in_dis out_h out_h_n rst_h set_h vcc_io 
+ vgnd vpwr
*.PININFO hld_h_n:I in:I in_dis:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr:I 
*.PININFO out_h:O out_h_n:O
XI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI34 in_i in_i_n virt_pwr vpwr sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 in_i_n in virt_pwr vpwr sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 virt_pwr in_dis vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI33 virt_pwr in_dis vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 in_i_n in_dis vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 in_i in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI58 net153 vpwr net113 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI59 net145 vpwr net117 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 fbk_n hld_h_n net145 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 in_i_n in vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 in_i in_dis vgnd vgnd sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 fbk hld_h_n net153 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 net117 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 net113 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_ctl_hld enable_h hld_h_n hld_i_h_n hld_i_ovr_h hld_i_vpwr 
+ hld_ovr od_i_h vcc_io vgnd vpwr
*.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h_n:O 
*.PININFO hld_i_ovr_h:O hld_i_vpwr:O od_i_h:O
Xhld_i_h_inv8<1> hld_i_h hld_i_h_n vgnd vgnd vcc_io vcc_io
+ sky130_fd_io__sio_hvsbt_inv_x8
Xhld_i_h_inv8<0> hld_i_h hld_i_h_n vgnd vgnd vcc_io vcc_io
+ sky130_fd_io__sio_hvsbt_inv_x8
Xhld_i_h_inv4 hld_i_h_n_ls hld_i_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x4
XI33 od_i_h_n od_i_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x4
XI36 od_h enable_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI35 od_h enable_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xhld_i_vpwr_inv hld_i_vpwr_n hld_i_vpwr vgnd vgnd vpwr vpwr 
+ sky130_fd_io__sio_lvlp_inv_x4
XI30 od_i_h hld_i_ovr_h_n hld_i_ovr_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nor
XI26 hld_i_h_n_ls hld_ovr_h hld_i_ovr_h_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nor
Xhld_i_h_inv1 hld_i_h_ls hld_i_h_n_ls vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x1
XI31 od_h od_i_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
Xhld_nand enable_h hld_h_n hld_i_h_ls vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xhld_i_vpwr_ls hld_i_h_n_ls hld_i_h_ls hld_i_vpwr_n net91 vgnd vpwr 
+ sky130_fd_io__sio_ctl_ls_out
Xanalog_en_ls hld_i_h_n_ls hld_ovr vgnd hld_ovr_h net101 vgnd vgnd vcc_io vgnd 
+ vpwr sky130_fd_io__sio_ctl_ls
.ENDS

.SUBCKT sky130_fd_io__sio_tk_opto out spd spu
*.PININFO out:B spd:B spu:B
Xe1 spu out sky130_fd_io__sio_tk_em1o
Xe2 out spd sky130_fd_io__sio_tk_em1s
.ENDS

.SUBCKT sky130_fd_io__sio_tk_opti out spd spu
*.PININFO out:B spd:B spu:B
Xe1 out spu sky130_fd_io__sio_tk_em1s
Xe2 spd out sky130_fd_io__sio_tk_em1o
.ENDS

.SUBCKT sky130_fd_io__sio_tk_optiA out spd spu
*.PININFO out:B spd:B spu:B
Xe1 out spu sky130_fd_io__sio_tk_em2s
Xe2 spd out sky130_fd_io__sio_tk_em1o
.ENDS

.SUBCKT sky130_fd_io__sio_ctl_lsbank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n hld_i_vpwr ibuf_sel ibuf_sel_h 
+ ibuf_sel_h_n inp_dis inp_dis_h inp_dis_h_n od_i_h vcc_io vgnd vpwr vtrip_sel 
+ vtrip_sel_h vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I hld_i_h_n:I hld_i_vpwr:I ibuf_sel:I 
*.PININFO inp_dis:I od_i_h:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I dm_h<2>:O 
*.PININFO dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O ibuf_sel_h:O 
*.PININFO ibuf_sel_h_n:O inp_dis_h:O inp_dis_h_n:O vtrip_sel_h:O 
*.PININFO vtrip_sel_h_n:O
Xdm_ls<2> hld_i_h_n dm<2> hld_i_vpwr dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> 
+ vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls
Xdm_ls<1> hld_i_h_n dm<1> hld_i_vpwr dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> 
+ vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls
Xdm_ls<0> hld_i_h_n dm<0> hld_i_vpwr dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> 
+ vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls
Xinp_dis_ls net81 inp_dis hld_i_vpwr inp_dis_h inp_dis_h_n ie_n_rst_h 
+ ie_n_st_h vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls
Xbuf_sel_ls hld_i_h_n ibuf_sel hld_i_vpwr ibuf_sel_h ibuf_sel_h_n 
+ buf_sel_rst_h buf_sel_st_h vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls
Xtrip_sel_ls hld_i_h_n vtrip_sel hld_i_vpwr vtrip_sel_h vtrip_sel_h_n 
+ trip_sel_rst_h trip_sel_st_h vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls

XI101 net81 hld_i_h_n vcc_io sky130_fd_io__sio_tk_opto
Xtrip_sel_st trip_sel_st_h od_i_h vgnd sky130_fd_io__sio_tk_opti
Xbuf_sel_rst buf_sel_rst_h vgnd od_i_h sky130_fd_io__sio_tk_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h sky130_fd_io__sio_tk_opti
Xdm_rst<2> dm_rst_h<2> vgnd od_i_h sky130_fd_io__sio_tk_opti
Xie_n_rst ie_n_rst_h vgnd od_i_h sky130_fd_io__sio_tk_opti
XI345<1> dm_st_h<1> od_i_h vgnd sky130_fd_io__sio_tk_opti
Xbuf_sel_st buf_sel_st_h od_i_h vgnd sky130_fd_io__sio_tk_opti
Xie_n_st ie_n_st_h od_i_h vgnd sky130_fd_io__sio_tk_opti
XI347<1> dm_rst_h<0> vgnd od_i_h sky130_fd_io__sio_tk_opti
Xdm_rst<1> dm_rst_h<1> vgnd od_i_h sky130_fd_io__sio_tk_opti
XI344<1> dm_st_h<0> od_i_h vgnd sky130_fd_io__sio_tk_opti
XI346<1> dm_st_h<2> od_i_h vgnd sky130_fd_io__sio_tk_opti

.ENDS

.SUBCKT sky130_fd_io__sio_ctl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> 
+ dm_h_n<1> dm_h_n<0> enable_h hld_h_n hld_i_h_n hld_i_ovr_h hld_i_vpwr 
+ hld_ovr ibuf_sel ibuf_sel_h ibuf_sel_h_n inp_dis inp_dis_h inp_dis_h_n 
+ od_i_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I hld_h_n:I hld_ovr:I ibuf_sel:I 
*.PININFO inp_dis:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I dm_h<2>:O dm_h<1>:O 
*.PININFO dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O hld_i_h_n:O 
*.PININFO hld_i_ovr_h:O hld_i_vpwr:O ibuf_sel_h:O ibuf_sel_h_n:O inp_dis_h:O 
*.PININFO inp_dis_h_n:O od_i_h:O vtrip_sel_h:O vtrip_sel_h_n:O
Xhld_dis_blk enable_h hld_h_n hld_i_h_n hld_i_ovr_h hld_i_vpwr hld_ovr od_i_h 
+ vcc_io vgnd vpwr sky130_fd_io__sio_ctl_hld
Xls_bank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hld_i_vpwr ibuf_sel ibuf_sel_h ibuf_sel_h_n inp_dis 
+ inp_dis_h inp_dis_h_n od_i_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h 
+ vtrip_sel_h_n sky130_fd_io__sio_ctl_lsbank
.ENDS

.SUBCKT sky130_fd_io__sio_pupredrvr_reg drvhi_h pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XI3 pu_h_n drvhi_h net27 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI39 net27 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pupredrvr_reg_slow drvhi_h pu_h_n puen_h slow_h_n vcc_io 
+ vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n:O
XI3 pu_h_n drvhi_h net34 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI39 net34 puen_h net30 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI61 net30 slow_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI60 pu_h_n slow_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_obpredrvr_reg drvhi_h pu_h_n<5> pu_h_n<4> puen_h slow_h_n 
+ vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<5>:O 
*.PININFO pu_h_n<4>:O
Xpu_reg drvhi_h pu_h_n<5> puen_h vcc_io vgnd_io sky130_fd_io__sio_pupredrvr_reg
XI73 drvhi_h pu_h_n<4> puen_h slow_h_n vcc_io vgnd_io 
+ sky130_fd_io__sio_pupredrvr_reg_slow
.ENDS

.SUBCKT sky130_fd_io__sio_com_pdpredrvr_pbias drvlo_h_n en_h en_h_n pbias pd_h 
+ pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_h:I en_h_n:I pd_h:I pden_h_n:I vcc_io:I vgnd_io:I 
*.PININFO pbias:O
XI27 n<0> pd_h en_h_n sky130_fd_io__sio_tk_opto
XE1 n<1> n<0> sky130_fd_io__sio_tk_em1o
XE2 pbias pbias1 sky130_fd_io__sio_tk_em1o
XE3 pbias1 net97 sky130_fd_io__sio_tk_em1s
XE4 net112 pbias sky130_fd_io__sio_tk_em1s
XE6 pbias net93 sky130_fd_io__sio_tk_em1s
XE5 n<101> bias_g sky130_fd_io__sio_tk_em1s
XI47 pbias bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 n<1> drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI18 bias_g drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI23 n<0> n<0> n<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 drvlo_i_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI20 bias_g n<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI19 bias_g en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI34 net169 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI36 net112 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI38 n<1> pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI48 n<100> pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI41 n<101> pd_h n<100> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI44 pbias pbias pbias1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI45 pbias1 pbias1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI15 net195 en_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI16 net183 n<0> net195 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 pbias en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 drvlo_i_h drvlo_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 bias_g drvlo_h_n net183 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI14 pbias drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI33 N0 vgnd_io vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 net173 net173 N0 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 net169 net169 net173 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 net97 N0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI43 net93 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI40 N0 drvlo_i_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
Xmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin_fast<1> pd_h drvlo_h_n int_nor<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin_fast<0> pd_h drvlo_h_n int_nor<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pdpredrvr_strong_nr2_i2c drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
Xmpin_slow pd_h drvlo_h_n int_slow vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_slow int_slow pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin_fast<1> pd_h drvlo_h_n int_nor<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin_fast<0> pd_h drvlo_h_n int_nor<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_inv_x1_dnw in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XI1 out in vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 out in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_nor2_dnw in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XI3 net17 in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out in1 net17 vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 out in1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pdpredrvr_strong drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> 
+ pd_h<2> pden_h_n slow_h vcc_io vgnd_io
*.PININFO drvlo_h_n:I i2c_mode_h_n:I pden_h_n:I slow_h:I vcc_io:I vgnd_io:I 
*.PININFO pd_h<4>:O pd_h<3>:O pd_h<2>:O
Xbias drvlo_h_n en_fast_h net167 pbias1 pd_h<2> pden_h_n vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pdpredrvr_pbias
Xnr2 drvlo_h_n en_fast2_n<1> en_fast2_n<0> pd_h<3> pden_h_n vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pdpredrvr_strong_nr2
Xnr3 drvlo_h_n net179 net179 pd_h<2> pden_h_n vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pdpredrvr_strong_nr2
XI93 net126 en_fast5_n<1> en_fast5_n<0> pd_h<4> i2c_mode_enable_h_n vcc_io 
+ vgnd_io sky130_fd_io__sio_com_pdpredrvr_strong_nr2_i2c
XI1 net128 i2c_mode_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net128 pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI118 net126 net136 vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI128 i2c_mode_enable_h_n net128 vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI117 net136 drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI3 net147 i2c_mode_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI130 net128 pden_h_n net147 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI119 net126 net136 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI129 i2c_mode_enable_h_n net128 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI115 net136 drvlo_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xinv en_fast_h net167 vgnd_io vcc_io sky130_fd_io__sio_com_inv_x1_dnw
XI86 slow_h pden_h_n en_fast_h vgnd_io vcc_io sky130_fd_io__sio_com_nor2_dnw
XI77 en_fast2_n<1> pbias1 net167 sky130_fd_io__sio_tk_opto
XI76 net179 pbias1 net167 sky130_fd_io__sio_tk_opto
XI94 en_fast5_n<1> pbias1 net167 sky130_fd_io__sio_tk_opto
XI96 en_fast5_n<0> en_fast5_n<1> vcc_io sky130_fd_io__sio_tk_optiA
XI79 en_fast2_n<0> en_fast2_n<1> vcc_io sky130_fd_io__sio_tk_opti
.ENDS

.SUBCKT sky130_fd_io__sio_com_pupredrvr_weak drvhi_h pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XI3 pu_h_n drvhi_h net21 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI39 net21 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pdpredrvr_weak drvlo_h_n pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
XI26 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI25 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 net25 pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI23 pd_h drvlo_h_n net25 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pupredrvr_strong_slow drvhi_h pu_h_n puen_h vcc_io 
+ vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XI3 pu_h_n drvhi_h net17 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI39 net17 puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI38 pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI37 pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pdpredrvr_strong_slow drvlo_h_n pd_h pden_h_n vcc_io 
+ vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
XI26 pd_h pden_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI25 pd_h drvlo_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 net25 pden_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI23 pd_h drvlo_h_n net25 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pupredrvr_nbias drvhi_h en_h en_h_n nbias pu_h_n 
+ puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_h:I en_h_n:I pu_h_n:I puen_h:I vcc_io:I vgnd_io:I 
*.PININFO nbias:O
XI36 n<2> pu_h_n en_h sky130_fd_io__sio_tk_opto
XE1 n<2> n<1> sky130_fd_io__sio_tk_em1o
XE2 n<6> nbias sky130_fd_io__sio_tk_em1o
XE5 nbias net138 sky130_fd_io__sio_tk_em1s
XE4 n<6> net236 sky130_fd_io__sio_tk_em1s
XE7 bias_g net132 sky130_fd_io__sio_tk_em1s
XE6 net192 nbias sky130_fd_io__sio_tk_em1s
XI34 n<1> drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 n<1> n<2> n<2> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 bias_g n<1> vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 bias_g drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI29 bias_g en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI21 nbias bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 drvhi_i_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI47 n<7> bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI49 net138 bias_g vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI50 n<1> puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI56 vcc_io pu_h_n net132 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI19 n<6> n<6> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI20 nbias nbias n<6> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI28 bias_g drvhi_h n<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI27 n<3> n<2> n<4> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI26 n<4> en_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 drvhi_i_h_n drvhi_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI24 nbias en_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI53 vccio_2vtn drvhi_i_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI25 nbias drvhi_i_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI40 vccio_2vtn vcc_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI39 net236 vccio_2vtn vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI44 n<8> n<8> vccio_2vtn vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI41 n<7> n<7> n<8> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI54 net192 bias_g vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XE1 net024 pu_h_n sky130_fd_io__sio_tk_em1s
XRrespu1 int_res net024 sky130_fd_pr__res_generic_po m=1 w=0.33 l=11
XRrespu2 pu_h_n int_res sky130_fd_pr__res_generic_po m=1 w=0.33 l=4
Xmnin_fast<3> net024 drvhi_h int<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_fast<2> net024 drvhi_h int<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_fast<1> net024 drvhi_h int<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_fast<0> net024 drvhi_h int<0> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_slow1 n<2> puen_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnin_slow pu_h_n drvhi_h n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<3> int<3> en_fast<3> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<2> int<2> en_fast<2> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<1> int<1> en_fast<1> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpen pu_h_n puen_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmpin pu_h_n drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_nand2_dnw in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XI3 out in0 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 out in1 vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in1 net25 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 net25 in0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h 
+ slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O
Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pupredrvr_nbias
Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> 
+ pu_h_n<3> puen_h vcc_io vgnd_io sky130_fd_io__sio_com_pupredrvr_strong_nd2
Xnd2a drvhi_h net57 net57 net57 net57 pu_h_n<2> puen_h vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pupredrvr_strong_nd2
XI102 puen_h slow_h_n en_fast_h_n vgnd_io vcc_io sky130_fd_io__sio_com_nand2_dnw
Xinv en_fast_h_n en_fast_h vgnd_io vcc_io sky130_fd_io__sio_com_inv_x1_dnw
XI92 en_fast_h_3<3> nbias_out en_fast_h sky130_fd_io__sio_tk_opto
XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io sky130_fd_io__sio_tk_opto
XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io sky130_fd_io__sio_tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io sky130_fd_io__sio_tk_opto
XI93 net57 nbias_out en_fast_h sky130_fd_io__sio_tk_opto
.ENDS

.SUBCKT sky130_fd_io__sio_obpredrvr drvhi_h drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> slow_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I i2c_mode_h_n:I pden_h_n<1>:I pden_h_n<0>:I 
*.PININFO puen_h<1>:I puen_h<0>:I slow_h:I slow_h_n:I vcc_io:I vgnd_io:I 
*.PININFO pd_h<4>:O pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O
Xpd_strong drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> pd_h<2> pden_h_n<1> slow_h 
+ vcc_io vgnd_io sky130_fd_io__sio_pdpredrvr_strong
Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pupredrvr_weak
Xpd_weak drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pdpredrvr_weak
Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pupredrvr_strong_slow
Xpd_strong_slow drvlo_h_n pd_h<1> pden_h_n<1> vcc_io vgnd_io 
+ sky130_fd_io__sio_com_pdpredrvr_strong_slow
Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io 
+ sky130_fd_io__sio_pupredrvr_strong
.ENDS

.SUBCKT sky130_fd_io__sio_hvsbt_xor in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XI3 net31 in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 out net56 net47 vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI17 net72 in1 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI18 net56 in0 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 net47 in1 vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out net72 net31 vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 out in1 net60 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI16 net72 in1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 out net72 net64 vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI15 net64 net56 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI14 net60 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI19 net56 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_octl_tsg4 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hld_i_vpwr od_h pden_h_n<2> pden_h_n<1> pden_h_n<0> 
+ puen_0_h puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd 
+ vpwr vreg_en_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_vpwr:I od_h:I slow:I vcc_io:I vgnd:I vpwr:I 
*.PININFO vreg_en_h_n:I pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O 
*.PININFO puen_2or1_h:O puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O
XI210 dm_h<2> dm_h<0> n<8> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_xor
XI200 dm_h<2> dm_h<1> n<10> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_xor
XI209 n<5> n<2> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI344 pden_h_n<2> net241 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI254 puen_h1_n puen_h<1> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI256 puen_h0_n puen_h<0> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI249 pden_h0 pden_h_n<0> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI247 pden_h1 pden_h_n<1> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI185 dm_h_n<0> n<4> net130 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI187 dm_h<1> dm_h<0> n<3> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI255 puen_0_h puen_0_h puen_h0_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI253 n<2> n<2> puen_h1_n vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI203 n<10> dm_h<0> n<1> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI204 n<9> dm_h_n<0> n<0> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI205 n<1> n<0> puen_2or1_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI365 net198 dm_h<2> pden_h_n<2> vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI211 n<8> dm_h_n<1> puen_0_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
XI246 net130 net130 pden_h1 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
XI248 n<3> n<3> pden_h0 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
XI366 dm_h<1> dm_h<0> net198 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
Xls_slow hld_i_h_n slow hld_i_vpwr slow_h slow_h_n od_h vgnd vcc_io vgnd vpwr 
+ sky130_fd_io__sio_ctl_ls
.ENDS

.SUBCKT sky130_fd_io__sio_octl_tsg4 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hld_i_vpwr od_h oe_h oe_hs_h pden_h_n<2> pden_h_n<1> 
+ pden_h_n<0> puen_h<2> puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd 
+ vpwr vreg_en vreg_en_h
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_vpwr:I od_h:I oe_h:I slow:I vcc_io:I vgnd:I vpwr:I 
*.PININFO vreg_en:I oe_hs_h:O pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O 
*.PININFO puen_h<2>:O puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O vreg_en_h:O
XI351 net125 puen_2or1_h n<1> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
XI352 n<1> oe_i_h_n oe_hs_i_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nor
XI353 oe_h oe_i_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI251 puen_h2_n puen_h<2> vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI355 oe_hs_i_h_n oe_hs_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x2
XI207 vreg_puen2 vreg_puen2_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x1
XI354 oe_hs_i_h oe_hs_i_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI206 puen_2or1_h vreg_en_h vreg_puen2 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI250 vreg_puen2_n vreg_puen2_n puen_h2_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
Xls_vreg_en hld_i_h_n vreg_en hld_i_vpwr vreg_en_h vreg_en_h_n od_h vgnd 
+ vcc_io vgnd vpwr sky130_fd_io__sio_ctl_ls
XI367 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_vpwr od_h pden_h_n<2> pden_h_n<1> pden_h_n<0> net125 puen_2or1_h 
+ puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd vpwr vreg_en_h_n 
+ sky130_fd_io__sio_com_octl_tsg4
.ENDS

.SUBCKT sky130_fd_io__sio_com_ls_nor2 in in_dis out vgnd virt_pwr vnb vpb vpwr
*.PININFO in:I in_dis:I vgnd:I vnb:I vpb:I vpwr:I out:O virt_pwr:B
Xnin out in vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xnen out in_dis vgnd vnb sky130_fd_pr__nfet_01v8 m=1 w=1.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpen virt_pwr in_dis vpwr vpb sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpin out in virt_pwr vpb sky130_fd_pr__pfet_01v8 m=1 w=3.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_dat_ls hld_h_n in in_dis out_h out_h_n rst_h set_h 
+ vcc_io vgnd vpwr_ka
*.PININFO hld_h_n:I in:I in_dis:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr_ka:I 
*.PININFO out_h:O out_h_n:O
Xnr1 in in_dis in_i_n vgnd virt_pwr vgnd vpwr_ka vpwr_ka 
+ sky130_fd_io__sio_com_ls_nor2
Xnr2 in_i_n in_dis in_i vgnd virt_pwr vgnd vpwr_ka vpwr_ka 
+ sky130_fd_io__sio_com_ls_nor2
XI3 fbk fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 fbk hld_h_n net81 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI6 fbk_n hld_h_n net85 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI7 net109 in_i_n vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=8 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI8 net105 in_i vgnd vgnd sky130_fd_pr__nfet_01v8_lvt m=8 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI12 out_h fbk_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI13 out_h_n fbk vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnset fbk_n set_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmnrst fbk rst_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI31 net85 vpwr_ka net105 vgnd sky130_fd_pr__nfet_05v0_nvt m=8 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI30 net81 vpwr_ka net109 vgnd sky130_fd_pr__nfet_05v0_nvt m=8 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI11 out_h fbk_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI14 out_h_n fbk vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_cclat_hvnand3 in0 in1 in2 out vcc_io vgnd vnb
*.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
Xmp0 out in0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmp2 out in2 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmp1 out in1 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmn2 out in2 n1 vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
Xmn0 n0 in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmn1 n1 in1 n0 vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_cclat_hvnor3 in0 in1 in2 out vcc_io vgnd vnb
*.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
Xmp0 n<0> in0 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmp2 out in2 n<1> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmp1 n<1> in1 n<0> vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmn0 out in0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmn2 out in2 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmn1 out in1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_cclat_inv_in in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
Xmp1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xmn1 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_cclat_inv_out in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XI1 out in vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=6 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI2 out in vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_cclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io 
+ vgnd
*.PININFO oe_h_n:I pd_dis_h:I pu_dis_h:I vcc_io:I vgnd:I drvhi_h:O drvlo_h_n:O
Xnand3 oe_i_h drvlo_h_n pu_dis_h_n n0 vcc_io vgnd vgnd 
+ sky130_fd_io__sio_com_cclat_hvnand3
Xnor3 oe_i_h_n drvhi_h pd_dis_h n1 vcc_io vgnd vgnd 
+ sky130_fd_io__sio_com_cclat_hvnor3
Xinv_oe1 oe_h_n oe_i_h vcc_io vgnd vgnd sky130_fd_io__sio_com_cclat_inv_in
Xinv_oe2 oe_i_h oe_i_h_n vcc_io vgnd vgnd sky130_fd_io__sio_com_cclat_inv_in
Xinv_pudis pu_dis_h pu_dis_h_n vcc_io vgnd vgnd sky130_fd_io__sio_com_cclat_inv_in
Xinv_out n1 drvlo_h_n vcc_io vgnd vgnd sky130_fd_io__sio_com_cclat_inv_out
Xinv_out_1 n0 drvhi_h vcc_io vgnd vgnd sky130_fd_io__sio_com_cclat_inv_out
.ENDS

.SUBCKT sky130_fd_io__sio_opath_datoe din drvhi_h drvlo_h_n hld_i_ovr_h od_h oe_h 
+ oe_n vcc_io vgnd vpwr_ka
*.PININFO din:I hld_i_ovr_h:I od_h:I oe_n:I vcc_io:I vgnd:I vpwr_ka:I 
*.PININFO drvhi_h:O drvlo_h_n:O oe_h:O
Xdat_ls hld_i_ovr_h din vgnd pd_dis_h pu_dis_h vgnd od_h vcc_io vgnd vpwr_ka 
+ sky130_fd_io__sio_com_dat_ls
Xoe_ls hld_i_ovr_h oe_n vgnd oe_h_n oe_h vgnd od_h vcc_io vgnd vpwr_ka 
+ sky130_fd_io__sio_com_dat_ls
Xcclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io vgnd 
+ sky130_fd_io__sio_cclat
.ENDS

.SUBCKT sky130_fd_io__sio_octl_dat din dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h hld_i_vpwr od_h oe_hs_h oe_n pd_h<4> 
+ pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> 
+ puen_h<2> slow slow_h_n vcc_io vgnd vgnd_io vpwr vpwr_ka vreg_en vreg_en_h
*.PININFO din:I dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I 
*.PININFO dm_h_n<0>:I hld_i_h_n:I hld_i_ovr_h:I hld_i_vpwr:I od_h:I oe_n:I 
*.PININFO slow:I vcc_io:I vgnd:I vgnd_io:I vpwr:I vpwr_ka:I vreg_en:I 
*.PININFO drvhi_h:O oe_hs_h:O pd_h<4>:O pd_h<3>:O pd_h<2>:O pd_h<1>:O 
*.PININFO pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O 
*.PININFO puen_h<2>:O slow_h_n:O vreg_en_h:O
Xpredrvr drvhi_h drvlo_h_n pden_h_n<2> pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
+ puen_h<0> slow_h slow_h_n vcc_io vgnd_io sky130_fd_io__sio_obpredrvr
Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_vpwr od_h oe_h oe_hs_h pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_h<2> 
+ puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd vpwr vreg_en vreg_en_h 
+ sky130_fd_io__sio_octl_tsg4
Xdatoe din drvhi_h drvlo_h_n hld_i_ovr_h od_h oe_h oe_n vcc_io vgnd vpwr_ka 
+ sky130_fd_io__sio_opath_datoe
.ENDS

.SUBCKT sky130_fd_io__sio_opath_sub din dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h hld_i_vpwr od_h oe_hs_h oe_n pd_h<4> 
+ pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<5> pu_h_n<4> pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_reg_h slow slow_h_n vcc_io vgnd vgnd_io vpwr 
+ vpwr_ka vreg_en vreg_en_h
*.PININFO din:I dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I 
*.PININFO dm_h_n<0>:I hld_i_h_n:I hld_i_ovr_h:I hld_i_vpwr:I od_h:I oe_n:I 
*.PININFO slow:I vcc_io:I vgnd:I vgnd_io:I vpwr:I vpwr_ka:I vreg_en:I 
*.PININFO drvhi_h:O oe_hs_h:O pd_h<4>:O pd_h<3>:O pd_h<2>:O pd_h<1>:O 
*.PININFO pd_h<0>:O pu_h_n<5>:O pu_h_n<4>:O pu_h_n<3>:O pu_h_n<2>:O 
*.PININFO pu_h_n<1>:O pu_h_n<0>:O puen_reg_h:O slow_h_n:O vreg_en_h:O
Xpredrvr_reg drvhi_h pu_h_n<5> pu_h_n<4> puen_reg_h slow_h_n vcc_io vgnd_io 
+ sky130_fd_io__sio_obpredrvr_reg
Xopath din dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h 
+ hld_i_h_n hld_i_ovr_h hld_i_vpwr od_h oe_hs_h oe_n pd_h<4> pd_h<3> pd_h<2> 
+ pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_reg_h slow 
+ slow_h_n vcc_io vgnd vgnd_io vpwr vpwr_ka vreg_en vreg_en_h 
+ sky130_fd_io__sio_octl_dat
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_nonoverlap p1g p2g padlo vgnd vpwr
*.PININFO padlo:I vgnd:I vpwr:I p1g:O p2g:O
XI76 p1g p1gb vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI64 p1g_new padlo vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI53 padlo_bar padlo vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI50 p2g_new p1g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI49 p2g_new padlo_bar vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI65 p1g_new p2g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI77 p2g p2gb vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI70 p2gb p2g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI72 p1gb p1g_new vpwr vpwr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI54 padlo_bar padlo vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI69 p1g_new padlo net140 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI78 p2g p2gb vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI67 net140 p2g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI71 p2gb p2g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI79 p1g p1gb vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI51 p2g_new padlo_bar net124 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI73 p1gb p1g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI52 net124 p1g_new vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_bias pswg_h vcc_io vpb_drvr
*.PININFO pswg_h:I vcc_io:I vpb_drvr:O
Xpsw_vccio vpb_drvr pswg_h vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=24 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_pug pad padlo pug_h tie_hi vpb_drvr
*.PININFO pad:I padlo:I tie_hi:I vpb_drvr:I pug_h:O
XEs1 pad net19 sky130_fd_io__tk_em1o
XEg2 net25 net21 sky130_fd_io__tk_em1o
XEg1 padlo net25 sky130_fd_io__tk_em1s
XI65 net21 tie_hi sky130_fd_io__tk_em1s
XEs2 net19 tie_hi sky130_fd_io__tk_em1s
XI52 pug_h net25 net19 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=1.825 sb=1.825 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI53 pug_h net21 net19 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_pghspu pad pghs_h pghs_h_latch tie_hi vcc_io_soft 
+ vpb_drvr
*.PININFO pad:I tie_hi:I vcc_io_soft:I vpb_drvr:I pghs_h:O pghs_h_latch:O
XEg9 tie_hi pg8 sky130_fd_io__tk_em1o
XEpghs6 pghs_h padhi6 sky130_fd_io__tk_em1s
XEg6 pg6 pg5 sky130_fd_io__tk_em1s
XEg2 pg2 pg1 sky130_fd_io__tk_em1s
XEg5 pg5 pg4 sky130_fd_io__tk_em1s
XEg4 pg4 pg3 sky130_fd_io__tk_em1s
XEpghs5 pghs_h padhi5 sky130_fd_io__tk_em1s
XEg1 pg1 vcc_io_soft sky130_fd_io__tk_em1s
XEpghs3 pghs_h_latch padhi3 sky130_fd_io__tk_em1s
XEg3 pg3 pg2 sky130_fd_io__tk_em1s
XEpghs7 pghs_h padhi7 sky130_fd_io__tk_em1s
XEg7 pg7 pg6 sky130_fd_io__tk_em1s
XEg8 pg8 pg7 sky130_fd_io__tk_em1s
XEpghs2 pghs_h_latch padhi2 sky130_fd_io__tk_em1s
XEpghs1 pghs_h_latch padhi1 sky130_fd_io__tk_em1s
XEpghs4 pghs_h_latch padhi4 sky130_fd_io__tk_em1s
XEpghs8 pghs_h padhi8 sky130_fd_io__tk_em1s
Xpghs5 padhi5 pg5 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs1 padhi1 pg1 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs8 padhi8 pg8 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs2 padhi2 pg2 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs3 padhi3 pg3 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs6 padhi6 pg6 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs4 padhi4 pg4 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpghs7 padhi7 pg7 pad vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_latch dishs_h dishs_h_n enhs_h enhs_h_n 
+ enhs_lat_h_n enhs_lathys_h_n exiths_h p3out pad_esd pghs_h vcc_io vgnd 
+ vpb_drvr vpwr_ka
*.PININFO dishs_h:I dishs_h_n:I enhs_h:I enhs_h_n:I exiths_h:I pad_esd:I 
*.PININFO vcc_io:I vgnd:I vpb_drvr:I vpwr_ka:I enhs_lat_h_n:O 
*.PININFO enhs_lathys_h_n:O p3out:O pghs_h:B
XI660 vgnd net102 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI528 n6 net96 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XEhys2 enhs_lathys_h_n enhs_lat_h_n sky130_fd_io__tk_em1o
XI658 net96 enhs_lat_h_n sky130_fd_io__tk_em1s
XEhys1 net117 enhs_lathys_h_n sky130_fd_io__tk_em1s
Xhys n6 net117 vcc_io vgnd sky130_fd_io__sio_hotswap_hys
Xpghspd enhs_h n2 pghs_h vgnd sky130_fd_io__sio_hotswap_pghspd
Xwpdenhs vpwr_ka net127 vgnd sky130_fd_io__sio_hotswap_wpd
Xwpdexhs vpwr_ka net124 vgnd sky130_fd_io__sio_hotswap_wpd
XI502 net186 pghs_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI484 net161 enhs_h pghs_h vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI491 n5 n6 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI498 n2 n6 net124 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI500 net170 enhs_h_n n2 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xnexiths pghs_h exiths_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI485 n3 n2 net161 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI499 n4 pghs_h net170 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI497 n6 n5 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xndishs pghs_h dishs_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI508 n2 enhs_h_n net186 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI696 vgnd exiths_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI487 pghs_h n5 net127 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI697 vgnd dishs_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI492 n5 n6 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI503 n4 vgnd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI488 n3 vgnd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI505 n6 n5 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI493 n5 n3 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI323 n2 dishs_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI279 n2 pad_esd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI504 n6 n4 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI689 p3out pad_esd vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=8 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_log dishs_h dishs_h_n en_h enhs_h enhs_h_n 
+ enhs_lat_h_n exiths_h forcehi_h<1> od_h vcc_io vgnd
*.PININFO en_h:I enhs_lat_h_n:I forcehi_h<1>:I od_h:I vcc_io:I vgnd:I 
*.PININFO dishs_h:O dishs_h_n:O enhs_h:O enhs_h_n:O exiths_h:O
XI664 net39 net46 dishs_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI663 od_h forcehi_h<1> net46 vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nand2
XI662 net62 en_h net39 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_nand2
XI658 od_h net62 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI666 enhs_lat_h_n net56 vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI565 net56 enhs_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI667 dishs_h dishs_h_n vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI637 enhs_h_n enhs_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
XI553 net56 enhs_dly_h_n exiths_h vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_nor
XI521 net56 enhs_dly_h enhs_dly_h_n vcc_io vgnd sky130_fd_io__sio_hotswap_dly
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_ctl en_h enhs_lat_h_n forcehi_h<1> od_h p3out 
+ pad_esd pghs_h vcc_io vgnd vpb_drvr vpwr_ka
*.PININFO en_h:I forcehi_h<1>:I od_h:I pad_esd:I vcc_io:I vgnd:I vpb_drvr:I 
*.PININFO vpwr_ka:I enhs_lat_h_n:O p3out:O pghs_h:B
Xhslatch dishs_h dishs_h_n enhs_h enhs_h_n enhs_lat_h_n enhs_lathys_h_n 
+ exiths_h p3out pad_esd pghs_h vcc_io vgnd vpb_drvr vpwr_ka 
+ sky130_fd_io__sio_hotswap_latch
Xhslog dishs_h dishs_h_n en_h enhs_h enhs_h_n enhs_lathys_h_n exiths_h 
+ forcehi_h<1> od_h vcc_io vgnd sky130_fd_io__sio_hotswap_log
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_pghs en_h force_h<1> od_h p3out pad padlo pghs_h 
+ tie_hi vcc_io vcc_io_soft vgnd vpb_drvr vpwr_ka
*.PININFO en_h:I force_h<1>:I od_h:I pad:I tie_hi:I vcc_io:I vcc_io_soft:I 
*.PININFO vgnd:I vpb_drvr:I vpwr_ka:I p3out:O padlo:O pghs_h:O
XI2 enhs_lat_h enhs_latbuf_h_n vgnd vgnd vcc_io vcc_io 
+ sky130_fd_io__sio_hvsbt_inv_x4
XI3 enhs_latbuf_h_n padlo sky130_fd_io__tk_em1s
XEpghs12 pghs_h net50 sky130_fd_io__tk_em1o
XI1 enhs_lat_h_n enhs_lat_h vgnd vgnd vcc_io vcc_io sky130_fd_io__sio_hvsbt_inv_x1
Xpghspu pad pghs_h net71 tie_hi vcc_io_soft vpb_drvr 
+ sky130_fd_io__sio_hotswap_pghspu
Xhsctl en_h enhs_lat_h_n force_h<1> od_h p3out pad net71 vcc_io vgnd vpb_drvr 
+ vpwr_ka sky130_fd_io__sio_hotswap_ctl
* Xclamp vgnd vcc_io vgnd vcc_io pad vgnd sky130_fd_io__signal_5_sym_hv_local_5term
Xclamp vgnd vcc_io vgnd vgnd pad vgnd sky130_fd_io__signal_5_sym_hv_local_5term
Xpghs12 net50 padlo vpb_drvr vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__res75only_noshorts_nometal pad rout
*.PININFO pad:B rout:B
XRI175 pad rout sky130_fd_pr__res_generic_po m=1 w=4 l=6.06
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap force_h<1> od_h oe_hs_h p2g pad pghs_h pug_h<5> 
+ pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> vcc_io vcc_io_soft vgnd 
+ vpb_drvr vpwr_ka
*.PININFO force_h<1>:I od_h:I oe_hs_h:I pad:I vcc_io:I vgnd:I vpwr_ka:I p2g:O 
*.PININFO pghs_h:O pug_h<5>:O pug_h<4>:O pug_h<3>:O pug_h<2>:O pug_h<1>:O 
*.PININFO pug_h<0>:O vcc_io_soft:O vpb_drvr:O
XI36 p1g p2g padlo vgnd vpb_drvr sky130_fd_io__sio_hotswap_nonoverlap
Xresd_tiehi vpb_drvr tie_hi sky130_fd_io__tk_tie_r_out_esd
Xresd_vccio vcc_io vcc_io_soft sky130_fd_io__tk_tie_r_out_esd
Xbias p1g vcc_io vpb_drvr sky130_fd_io__sio_hotswap_bias
Xpug<5> net102 net126 pug_h<5> tie_hi vpb_drvr sky130_fd_io__sio_hotswap_pug
Xpug<4> net102 net126 pug_h<4> tie_hi vpb_drvr sky130_fd_io__sio_hotswap_pug
Xpug<3> net102 net126 pug_h<3> tie_hi vpb_drvr sky130_fd_io__sio_hotswap_pug
Xpug<2> net102 net126 pug_h<2> tie_hi vpb_drvr sky130_fd_io__sio_hotswap_pug
Xpug<1> net102 net126 pug_h<1> tie_hi vpb_drvr sky130_fd_io__sio_hotswap_pug
Xpug<0> net102 net126 pug_h<0> tie_hi vpb_drvr sky130_fd_io__sio_hotswap_pug
Xpghs oe_hs_h force_h<1> od_h net95 net102 padlo net123 tie_hi vcc_io 
+ vcc_io_soft vgnd vpb_drvr vpwr_ka sky130_fd_io__sio_hotswap_pghs
XI113 pad net102 sky130_fd_io__res75only_noshorts_nometal
RI25 p1g net123 sky130_fd_pr__res_generic_m2 l=0.01 w=0.5
RI26 p2g net117 sky130_fd_pr__res_generic_m2 l=0.01 w=0.5
RI39 p2g net95 sky130_fd_pr__res_generic_m2 l=0.01 w=0.5
RI27 padlo net126 sky130_fd_pr__res_generic_m2 l=0.01 w=0.5
RI225 pghs_h p1g sky130_fd_pr__res_generic_m2 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__sio_tk_tie_r300 a b
*.PININFO a:B b:B
XRr1 a b sky130_fd_pr__res_generic_po m=1 w=0.5 l=3
.ENDS

.SUBCKT sky130_fd_io__sio_tk_tie_r a b
*.PININFO a:B b:B
Xres a b sky130_fd_io__sio_tk_tie_r300
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_unit pb pd pgin ps
*.PININFO pb:I pgin:I pd:B ps:B
Xpdrv pd pgin ps pb sky130_fd_pr__esd_pfet_g5v0d10v5 m=1 w=15.50 l=0.55 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_hotswap_vpb_bias p2g pad soft_vcc_io tie_hi vpb_drvr
*.PININFO p2g:I pad:I soft_vcc_io:I tie_hi:I vpb_drvr:B
XEpghs4 vpb_drvr net62 sky130_fd_io__tk_em1s
XEg3 net33 net37 sky130_fd_io__tk_em1s
XEpghs2 vpb_drvr net54 sky130_fd_io__tk_em1s
XEg4 net29 net33 sky130_fd_io__tk_em1s
XEg2 net37 net31 sky130_fd_io__tk_em1s
XEg5 net68 net29 sky130_fd_io__tk_em1s
XEpghs3 vpb_drvr net66 sky130_fd_io__tk_em1s
XEg1 p2g net31 sky130_fd_io__tk_em1s
XI5 tie_hi soft_vcc_io sky130_fd_io__tk_em1o
Xpsw_pad4 vpb_drvr net66 net68 pad sky130_fd_io__sio_pudrvr_unit
Xpsw_pad0 vpb_drvr net62 net31 pad sky130_fd_io__sio_pudrvr_unit
Xpsw_pad3 vpb_drvr net66 net29 pad sky130_fd_io__sio_pudrvr_unit
Xpsw_pad2 vpb_drvr net54 net33 pad sky130_fd_io__sio_pudrvr_unit
Xpsw_pad5 vpb_drvr vpb_drvr soft_vcc_io pad sky130_fd_io__sio_pudrvr_unit
Xpsw_pad1 vpb_drvr net54 net37 pad sky130_fd_io__sio_pudrvr_unit
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_strong_4 pad pug<3> pug<2> vcc_io vpb_drvr
*.PININFO vcc_io:I vpb_drvr:I pad:O pug<3>:B pug<2>:B
Xp5 vpb_drvr pad p5g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp6 vpb_drvr pad p6g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp7 vpb_drvr pad p7g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp8 vpb_drvr pad p8g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp4 vpb_drvr pad p4g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp3 vpb_drvr pad p3g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp2 vpb_drvr pad p2g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp1 vpb_drvr pad p1g vcc_io sky130_fd_io__sio_pudrvr_unit
XI35 p3g pug<3> pug<2> sky130_fd_io__sio_tk_opti
XI36 p4g pug<3> pug<2> sky130_fd_io__sio_tk_opti
XI33 p1g pug<3> pug<2> sky130_fd_io__sio_tk_opti
XI34 p2g pug<3> pug<2> sky130_fd_io__sio_tk_opti
XI42 p6g pug<3> pug<2> sky130_fd_io__sio_tk_opti
XI41 p5g pug<3> pug<2> sky130_fd_io__sio_tk_opti
XI44 p8g pug<3> pug<2> sky130_fd_io__sio_tk_opto
XI43 p7g pug<3> pug<2> sky130_fd_io__sio_tk_opto
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_strong nghs_h<3> nghs_h<2> p2gate pad pghs_h<3> 
+ pghs_h<2> pu_h_n<3> pu_h_n<2> pug<3> pug<2> vcc_io vcc_io_soft vgnd vgnd_io 
+ vpb_drvr
*.PININFO nghs_h<3>:I nghs_h<2>:I p2gate:I pghs_h<3>:I pghs_h<2>:I pu_h_n<3>:I 
*.PININFO pu_h_n<2>:I vcc_io:I vcc_io_soft:I vgnd:I vgnd_io:I vpb_drvr:I pad:O 
*.PININFO pug<3>:B pug<2>:B
XI190 p2gate pad vcc_io_soft tie_hi vpb_drvr sky130_fd_io__sio_hotswap_vpb_bias
XE6 p7g p6g sky130_fd_io__tk_em1o
XE11 p10g p11g sky130_fd_io__tk_em1o
XE4 p5g p4g sky130_fd_io__tk_em1s
XE13 p12g p13g sky130_fd_io__tk_em1s
XE3 p4g p3g sky130_fd_io__tk_em1s
XE12 p11g p12g sky130_fd_io__tk_em1s
XE1 p2g pug<2> sky130_fd_io__tk_em1s
XE2 p3g p2g sky130_fd_io__tk_em1s
XE14 p13g p14g sky130_fd_io__tk_em1s
XE10 p9g p10g sky130_fd_io__tk_em1s
XE20 tie_hi tie_hi_opt sky130_fd_io__tk_em1s
XE19 tie_hi p7g sky130_fd_io__tk_em1s
XE17 tie_hi_opt p17g sky130_fd_io__tk_em1s
XE8 p17g p8g sky130_fd_io__tk_em1s
XE9 tie_hi_opt p9g sky130_fd_io__tk_em1s
XE7 p8g p7g sky130_fd_io__tk_em1s
XE15 p14g p15g sky130_fd_io__tk_em1s
XE5 p6g p5g sky130_fd_io__tk_em1s
XE16 p15g pug<3> sky130_fd_io__tk_em1s
Xresd vpb_drvr tie_hi sky130_fd_io__sio_tk_tie_r_out_esd
Xp19 pad pug<3> pug<2> vcc_io vpb_drvr sky130_fd_io__sio_pudrvr_strong_4
Xp3 vpb_drvr pad p3g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp12 vpb_drvr pad p12g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp1 vpb_drvr pad pug<2> vcc_io sky130_fd_io__sio_pudrvr_unit
Xp2 vpb_drvr pad p2g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp4 vpb_drvr pad p4g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp18 vpb_drvr pad tie_hi vpb_drvr sky130_fd_io__sio_pudrvr_unit
Xp5 vpb_drvr pad p5g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp6 vpb_drvr pad p6g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp7 vpb_drvr pad p7g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp10 vpb_drvr pad p10g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp16 vpb_drvr pad pug<3> vcc_io sky130_fd_io__sio_pudrvr_unit
Xp15 vpb_drvr pad p15g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp14 vpb_drvr pad p14g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp9 vpb_drvr pad p9g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp8 vpb_drvr pad p8g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp13 vpb_drvr pad p13g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp11 vpb_drvr pad p11g vcc_io sky130_fd_io__sio_pudrvr_unit
Xp17 vpb_drvr pad p17g vcc_io sky130_fd_io__sio_pudrvr_unit
XI183 pug<3> nghs_h<3> pu_h_n<3> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI49 pug<2> nghs_h<2> pu_h_n<2> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI184 pu_h_n<3> pghs_h<3> pug<3> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI48 pu_h_n<2> pghs_h<2> pug<2> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_com_res_strong_slow ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
XE1 ra rb sky130_fd_io__sio_tk_em1o
XRr1 rb ra sky130_fd_pr__res_generic_po m=1 w=2 l=10
.ENDS

.SUBCKT sky130_fd_io__sio_pddrvr_unit nd ngin ns
*.PININFO ngin:I nd:B ns:B
Xndrv nd ngin ns ns sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=50.99 l=0.55 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pddrvr_strong pad pd_h<4> pd_h<3> pd_h<2> tie_lo_esd 
+ vcc_io vgnd_io
*.PININFO pd_h<4>:I pd_h<3>:I pd_h<2>:I vcc_io:I vgnd_io:I pad:O tie_lo_esd:O
XE9 tie_lo_esd ng<4> sky130_fd_io__tk_em2o
XE7 pd_h<4> ng<6> sky130_fd_io__tk_em1o
XE2 ng<2> ng<3> sky130_fd_io__tk_em1o
XE8 tie_lo_esd ng<3> sky130_fd_io__tk_em2o
XE6 tie_lo_esd ng<6> sky130_fd_io__tk_em2s
XE4 ng<4> pd_h<3> sky130_fd_io__tk_em1s
XE3 ng<3> ng<4> sky130_fd_io__tk_em1s
XE1 pd_h<2> ng<2> sky130_fd_io__tk_em1s
XI49 vgnd_io tie_lo_esd sky130_fd_io__sio_tk_tie_r_out_esd
Xn6 pad ng<6> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn5 pad pd_h<3> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn4 pad ng<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn3 pad ng<3> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn2 pad ng<2> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn1 pad pd_h<2> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<13> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<12> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<11> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<10> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<9> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<8> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<7> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<6> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<5> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<4> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<3> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<2> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<1> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
Xn8<0> pad pd_h<4> vgnd_io sky130_fd_io__sio_pddrvr_unit
RI8 vcc_io net76 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__sio_res_weak ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
Xe9 n<0> n<1> sky130_fd_io__sio_tk_em1s
Xe11 n<2> n<3> sky130_fd_io__sio_tk_em1s
Xe10 n<1> n<2> sky130_fd_io__sio_tk_em1s
Xe12 n<3> rb sky130_fd_io__sio_tk_em1s
Xe13 n<4> n<0> sky130_fd_io__sio_tk_em1s
Xe14 n<5> n<4> sky130_fd_io__sio_tk_em1o
XRI84 n<0> n<1> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
XRI62 n<3> rb sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
XRI82 n<2> n<3> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
XRI85 ra net64 sky130_fd_pr__res_generic_po m=1 w=0.8 l=50
XRI83 n<1> n<2> sky130_fd_pr__res_generic_po m=1 w=0.8 l=1.5
XRI116 net64 n<5> sky130_fd_pr__res_generic_po m=1 w=0.8 l=12
XRI104 n<4> n<0> sky130_fd_pr__res_generic_po m=1 w=0.8 l=6
XRI134 n<5> n<4> sky130_fd_pr__res_generic_po m=1 w=0.8 l=6
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_strong_slow pad pu_h_n vcc_io vgnd_io vpb_drvr
*.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
Xpdrv pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_weak pad pu_h_n vcc_io vgnd_io vpb_drvr
*.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
Xpdrv pad pu_h_n vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=8 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pddrvr_weak pad pd_h vcc_io vgnd_io
*.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
Xndrv1 pad pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pddrvr_strong_slow pad pd_h vcc_io vgnd_io
*.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
Xndrv pad pd_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_odrvr_nonreg nghs_h p2g pad pd_h<4> pd_h<3> pd_h<2> 
+ pd_h<1> pd_h<0> pghs_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug<3> pug<2> 
+ pug<1> pug<0> tie_lo_esd vcc_io vcc_io_soft vgnd vgnd_io vpb_drvr
*.PININFO nghs_h:I p2g:I pd_h<4>:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I 
*.PININFO pghs_h:I pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I 
*.PININFO vcc_io_soft:I vgnd:I vgnd_io:I vpb_drvr:I pad:O tie_lo_esd:O 
*.PININFO pug<3>:B pug<2>:B pug<1>:B pug<0>:B
Xpudrvr_strong nghs_h nghs_h p2g pad pghs_h pghs_h pu_h_n<3> pu_h_n<2> pug<3> 
+ pug<2> vcc_io vcc_io_soft vgnd vgnd_io vpb_drvr sky130_fd_io__sio_pudrvr_strong
Xresd pad_r250 pad sky130_fd_io__sio_res250only_small_esd
Xres pad_strong_slow pad_r250 vgnd_io sky130_fd_io__sio_com_res_strong_slow
Xpddrvr_strong pad pd_h<4> pd_h<3> pd_h<2> tie_lo_esd vcc_io vgnd_io 
+ sky130_fd_io__sio_pddrvr_strong
Xres_weak pad_weak pad_r250 vgnd_io sky130_fd_io__sio_res_weak
Xstrong_slow_pudrvr pad_strong_slow pug<1> vcc_io vgnd_io vpb_drvr 
+ sky130_fd_io__sio_pudrvr_strong_slow
Xpudrvr_weak pad_weak pug<0> vcc_io vgnd_io vpb_drvr sky130_fd_io__sio_pudrvr_weak
Xpddrvr_weak pad_weak pd_h<0> vcc_io vgnd_io sky130_fd_io__sio_pddrvr_weak
Xpddrvr pad_strong_slow pd_h<1> vcc_io vgnd_io 
+ sky130_fd_io__sio_pddrvr_strong_slow
XI50 pu_h_n<1> pghs_h pug<1> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI48 pu_h_n<0> pghs_h pug<0> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI51 pug<1> nghs_h pu_h_n<1> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI49 pug<0> nghs_h pu_h_n<0> vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_in_ctl_ls_out_reg in_c in_t out_c out_t vgnd vpb vpwr
*.PININFO in_c:I in_t:I vgnd:I vpb:I vpwr:I out_c:O out_t:O
XI35 out_c_n out_c vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 psa=265e-3 
+ pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 nw=1.00 nm=1
XI36 out_t_n out_t vgnd vgnd vpb vpwr sky130_fd_io__inv_p psd=280e-3 psb=265e-3 psa=265e-3 
+ pl=1.00 pw=1.00 pm=2 nsd=280e-3 nsb=265e-3 nsa=265e-3 nl=1.00 nw=1.00 nm=1
XI536 out_t_n in_t vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI535 out_c_n in_c vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.50 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI534 out_c_n out_t_n vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI533 out_t_n out_c_n vpwr vpb sky130_fd_pr__pfet_01v8 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__tk_em1o_b a b
*.PININFO a:B b:B
RI1 a net11 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI2 b net7 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__sio_tk_em1c a
*.PININFO a:B
RI1 a net10 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI2 a net6 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__sio_opamp_biasgen_reg ngate vgnd vpb vpwr vreg_en_n
*.PININFO vgnd:I vpb:I vpwr:I vreg_en_n:I ngate:B
XI201 net66 sky130_fd_io__sio_tk_em1c
XI206 net64 net70 sky130_fd_io__tk_em1o
XI235 net72 net64 sky130_fd_io__tk_em1o
XI234 net74 net72 sky130_fd_io__tk_em1o
XI207 net66 net74 sky130_fd_io__tk_em1o
XI208 ngate net66 sky130_fd_io__tk_em1o
XI187 net70 vreg_en_n vpwr vpb sky130_fd_pr__pfet_01v8 m=2 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> ngate ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> ngate ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xdummy vgnd vgnd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI334 ngate vreg_en_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XRI205 net66 net74 sky130_fd_pr__res_generic_po m=1 w=0.33 l=244.78
XRI199 net74 net72 sky130_fd_pr__res_generic_po m=1 w=0.33 l=282
XRR<0> net64 net70 sky130_fd_pr__res_generic_po m=1 w=0.33 l=253.63
XRI200 ngate net66 sky130_fd_pr__res_generic_po m=1 w=0.33 l=236.52
XRI203 net66 net66 sky130_fd_pr__res_generic_po m=1 w=0.33 l=47.06
XRI202 net72 net64 sky130_fd_pr__res_generic_po m=1 w=0.33 l=139.79
.ENDS

.SUBCKT sky130_fd_io__sio_opamp_stage_c_c_res b r1 r2
*.PININFO b:B r1:B r2:B
XI111 net36 r2 sky130_fd_io__sio_tk_em1s
XI474 net36 net41 sky130_fd_io__sio_tk_em1s
XI112 net40 net41 sky130_fd_io__sio_tk_em1o
XI113 net40 r1 sky130_fd_io__sio_tk_em1o
XRI91 net124 net76 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI54 r1 net49 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI89 net118 net109 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI88 net115 net124 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI55 net41 net46 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI90 net109 net52 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI86 net106 net118 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI98 net103 net36 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI97 net100 net36 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI110 net41 net88 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI109 r2 net91 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI108 net91 net82 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI107 net88 net85 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI106 net85 net73 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI105 net82 net79 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI104 net79 net67 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI92 net76 net58 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI103 net73 net70 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI102 net70 net61 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI101 net67 net64 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI100 net64 net100 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI99 net61 net103 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI95 net58 net40 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI94 net55 net40 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI93 net52 net55 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI85 net49 net106 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI84 net46 net43 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
XRI87 net43 net115 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=5
.ENDS

.SUBCKT sky130_fd_io__sio_opamp_stage_c_c en_hicc inn inp ngate out vcc vgnd vnb 
+ vpp vreg_en_h_n
*.PININFO en_hicc:I inn:I inp:I vcc:I vgnd:I vnb:I vpp:I vreg_en_h_n:I out:O 
*.PININFO ngate:B
XI491 vnb net_423 net_172 sky130_fd_io__sio_opamp_stage_c_c_res
XI456 vnb net400 out sky130_fd_io__sio_opamp_stage_c_c_res
XI490 vnb net356 net_172 sky130_fd_io__sio_opamp_stage_c_c_res
XI489 vnb net_339 out sky130_fd_io__sio_opamp_stage_c_c_res
XI472 net_435 pd_0 sky130_fd_io__tk_em1o
XI505 net315 vsource_1 sky130_fd_io__tk_em1o
XI470 pu_1 net_189 sky130_fd_io__tk_em1o
XI507 net327 vsource_0 sky130_fd_io__tk_em1o
XI468 net_391 pd_1 sky130_fd_io__tk_em1o
XI506 net315 vsource_1 sky130_fd_io__tk_em1o
XI475 pu_0 net_181 sky130_fd_io__tk_em1o
XI388 net_180 vsource_1 sky130_fd_io__tk_em1o
XI153 net_178 vsource_0 sky130_fd_io__tk_em1o
XI510 net327 vsource_0 sky130_fd_io__tk_em1o
XI444 vnb net315 sky130_fd_io__tk_em1s
XI509 vnb net327 sky130_fd_io__tk_em1s
XI473 vgnd net_435 sky130_fd_io__tk_em1s
XI471 net_189 net_233 sky130_fd_io__tk_em1s
XI474 net_181 vcc sky130_fd_io__tk_em1s
XI508 net327 vnb sky130_fd_io__tk_em1s
XI443 net315 vnb sky130_fd_io__tk_em1s
XI469 vgnd net_391 sky130_fd_io__tk_em1s
XI459 net_172 en_hicc_n out vpp sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<14> pd_0 net_307 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<12> net_307 net_307 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<13> pu_0 pu_0 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<8> out pu_0 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<9> out pu_0 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<10> out pu_0 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<11> out pu_0 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI360 net_172 en_hicc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI308 en_hicc_n en_hicc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI305 net_233 en_hicc_n vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI449 vcc net_181 vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<15> pd_1 net_444 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<17> net_444 net_444 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<16> pu_1 pu_1 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<18> net_172 pu_1 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<19> net_172 pu_1 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<20> net_172 pu_1 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<21> net_172 pu_1 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI266 net_233 net_189 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI463 vcc vcc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI462 net_233 net_233 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=3 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<25> net_307 vcc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<24> pu_0 vcc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI503 pd_0 vcc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI502 pd_1 net_233 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<23> net_444 net_233 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP1<22> pu_1 net_233 net_233 vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI511 pu_1 en_hicc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI513 net_444 en_hicc vcc vpp sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI460 out en_hicc net_172 vnb sky130_fd_pr__nfet_05v0_nvt m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<3> pu_0 inp vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<2> pu_0 inp vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<1> pu_0 inp vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<0> pu_0 inp vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI450 vgnd net_435 vgnd vnb sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<3> vsource_0 ngate vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI467 vgnd vgnd vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI415 pd_1 net_423 pd_1 pd_1 sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI413 net400 pu_0 net400 net400 sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<7> net_307 inn vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<6> net_307 inn vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<5> net_307 inn vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<4> net_307 inn vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI307 en_hicc_n en_hicc vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI466 net_398 vgnd vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<6> out pd_0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<7> out pd_0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<8> out pd_0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<9> out pd_0 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI492 net_398 vgnd vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<5> pd_0 pd_0 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI361 vgnd net_391 vgnd vnb sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI493 vgnd vgnd vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<11> pu_1 inp vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<10> pu_1 inp vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<9> pu_1 inp vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<8> pu_1 inp vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<4> vsource_1 ngate net_398 vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI422 net356 pu_1 net356 net356 sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<15> net_444 inn vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<14> net_444 inn vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<13> net_444 inn vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN1<12> net_444 inn vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI364 net_398 en_hicc vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<13> net_172 pd_1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<12> net_172 pd_1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<11> net_172 pd_1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<10> net_172 pd_1 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<14> pd_1 pd_1 vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM<7> net_180 ngate net_398 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<6> net_180 ngate net_398 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<5> net_180 ngate net_398 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI465 vsource_0 vsource_0 vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<2> net_178 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> net_178 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> net_178 ngate vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI464 vsource_0 vsource_0 vsource_0 net327 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI416 pd_0 net_339 pd_0 pd_0 sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI461 vsource_1 vsource_1 vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI458 vsource_1 vsource_1 vsource_1 net315 sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI501 out vreg_en_h_n vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI500 pd_1 en_hicc_n vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<15> pd_0 vgnd vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XMN<16> pd_1 vgnd vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_reg_opamp_c en_hicc fb_in fb_out refleak_bias 
+ vcc_io vgnd voutref vreg_en_h vreg_en_h_n
*.PININFO en_hicc:I fb_in:I refleak_bias:I vcc_io:I vgnd:I voutref:I 
*.PININFO vreg_en_h:I fb_out:O vreg_en_h_n:O
Xopamp_stage en_hicc fb_in voutref refleak_bias fb_out net30 vgnd vgnd vcc_io 
+ vreg_en_h_n sky130_fd_io__sio_opamp_stage_c_c
XI116 vreg_en_h_n vreg_en_h vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI117 net30 vreg_en_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI114 vreg_en_h_n vreg_en_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_reg_leak pad pu_h_n refleak_bias vcc_io vgnd_io
*.PININFO pu_h_n:I refleak_bias:I vcc_io:I vgnd_io:I pad:B
XE7 net35 net36 sky130_fd_io__tk_em1o
XE6 net31 net36 sky130_fd_io__tk_em1o
XI10 net51 net36 sky130_fd_io__tk_em1o
XE8 net75 net36 sky130_fd_io__tk_em1s
XE5 net37 net36 sky130_fd_io__tk_em1s
XI6 net55 pu_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xresd pad pad_esd sky130_fd_io__res250only_small
XML<14> net75 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<2> net37 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<1> net37 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<0> net37 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMEN pad_esd net55 net36 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<11> net31 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<10> net31 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<9> net31 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<8> net31 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<13> net35 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<12> net35 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI5 net55 pu_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XML<3> net51 refleak_bias vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xdummy vgnd_io vgnd_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_reg_csw_res b r1 r2
*.PININFO b:B r1:B r2:B
XI112 net40 net43 sky130_fd_io__tk_em1o
XI114 net40 r1 sky130_fd_io__tk_em1o
XI474 r2 net43 sky130_fd_io__tk_em1o
XRI126 net114 net45 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI54 r1 net48 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI89 net108 net102 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI125 net43 net63 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI90 net102 net51 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI130 net99 net96 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI129 net96 net69 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI86 net93 net108 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI121 net90 net84 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI124 net43 net72 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI123 net84 net81 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI122 net81 net75 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI120 net78 net66 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI119 net75 net78 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI118 net72 net90 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI132 net69 r2 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI117 net66 net40 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI131 net63 net54 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI115 net60 net40 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI94 net57 net60 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI128 net54 net114 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI93 net51 net57 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI85 net48 net93 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
XRI127 net45 net99 b sky130_fd_pr__res_generic_nd__hv m=1 w=0.33 l=4.4
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_reg_csw drvhi_h puen_reg_h slow_h_n vcc_io vgnd_io 
+ vpwr vref_nng vrefin
*.PININFO drvhi_h:I puen_reg_h:I slow_h_n:I vcc_io:I vgnd_io:I vpwr:I vrefin:I 
*.PININFO vref_nng:O
XI461 net214 vrefin sky130_fd_io__tk_em1o
XI387 vref_nng net76 sky130_fd_io__tk_em1o
XI395 net137 vrefin sky130_fd_io__tk_em1s
XI416 net125 vrefin sky130_fd_io__tk_em1s
XI396 vref_nng net82 sky130_fd_io__tk_em1s
XI417 vref_nng net80 sky130_fd_io__tk_em1s
XI418 vgnd_io int_5 nng_sd sky130_fd_io__sio_pudrvr_reg_csw_res
XI99 slow_h slow_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI284 psh_int_2 lvpsw_s psh_int_1 vpwr sky130_fd_pr__pfet_01v8 m=2 w=3.00 l=0.15 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI327 net82 hvpsw_s net137 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=8 w=3.00 l=0.50 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI385 puen_reg_h_n puen_reg_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI191 nng_sd drvhi_h_n_s vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI415 net80 hvpsw_s net125 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=16 w=3.00 l=0.50 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI368 hvpsw_s hvnsw_s vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI186 drvhi_h_n_s drvhi_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI280 hvnsw_s drvhi_h_n_s vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI324 drvhi_h_n_s puen_reg_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI414 int_5 slow_h_n nng_sd vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI380 int_1 slow_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI379 int_3 drvhi_h_n_s int_1 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI277 int_4 drvhi_h_n_s vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI378 int_3 vrefin vref_nng vgnd_io sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=2.00 mult=1 
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI374 ncap_s3 drvhi_h_n_s ncap_s2 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI290 vgnd_io ncap_s1 vgnd_io vgnd_io sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI281 hvnsw_s drvhi_h_n_s vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI190 int_5 vrefin vref_nng vgnd_io sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=2.00 mult=1 
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI100 slow_h slow_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI328 net214 hvnsw_s net76 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI367 hvpsw_s vpwr lvpsw_s vgnd_io sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI288 vgnd_io ncap_s2 vgnd_io vgnd_io sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI243 vrefin vpwr psh_int_1 vgnd_io sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI358 nng_sd drvhi_h_n_s int_4 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI187 drvhi_h_n_s drvhi_h int_2 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI326 psh_int_2 vpwr vref_nng vgnd_io sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI322 int_2 puen_reg_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI289 ncap_s3 ncap_s3 ncap_s2 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI293 vgnd_io ncap_s3 vgnd_io vgnd_io sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI295 vref_nng slow_h ncap_s3 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI369 hvpsw_s hvnsw_s vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=2 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI372 ncap_s2 drvhi_h_n_s vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI371 vref_nng slow_h ncap_s1 vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI386 puen_reg_h_n puen_reg_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI383 vref_nng puen_reg_h_n vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI370 ncap_s1 drvhi_h_n_s vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI430 lvpsw_s vgnd_io vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.00 l=0.50 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_esd_res pad rout
*.PININFO pad:B rout:B
XI2 pad rout sky130_fd_io__sio_tk_em1s
XRI175 pad rout sky130_fd_pr__res_generic_po m=1 w=2 l=10.41
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_reg_pu drvhi_h nghs_h pad pghs_h pu_h_n<1> 
+ pu_h_n<0> pug<1> pug<0> vcc_io vgnd vgnd_io vpb_drvr vref_int vref_nng
*.PININFO drvhi_h:I nghs_h:I pghs_h:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I vpb_drvr:I vref_int:I vref_nng:I pad:O pug<1>:B pug<0>:B
XI37 net134 vref_nng sky130_fd_io__tk_em1s
XI88 net196 net122 sky130_fd_io__tk_em1s
XI36 net249 net128 sky130_fd_io__tk_em1s
XI31 net132 vref_nng sky130_fd_io__tk_em1s
XI102 net221 net151 sky130_fd_io__tk_em1s
XI33<4> net253<0> net128 sky130_fd_io__tk_em1s
XI33<3> net253<1> net128 sky130_fd_io__tk_em1s
XI33<2> net253<2> net128 sky130_fd_io__tk_em1s
XI33<1> net253<3> net128 sky130_fd_io__tk_em1s
XI33<0> net253<4> net128 sky130_fd_io__tk_em1s
XI41 net144 net112 sky130_fd_io__tk_em1s
XI77 pad net110 sky130_fd_io__tk_em1s
XI99 net138 vref_nng sky130_fd_io__tk_em1s
XI84<1> net144 net106<0> sky130_fd_io__tk_em1s
XI84<0> net144 net106<1> sky130_fd_io__tk_em1s
XI97 net126 vref_nng sky130_fd_io__tk_em1s
XI106<3> net225<0> net128 sky130_fd_io__tk_em1s
XI106<2> net225<1> net128 sky130_fd_io__tk_em1s
XI106<1> net225<2> net128 sky130_fd_io__tk_em1s
XI106<0> net225<3> net128 sky130_fd_io__tk_em1s
XI89 net196 net140 sky130_fd_io__tk_em1o
XI100 net142 net138 sky130_fd_io__tk_em1o
XI43 net112 vref_nng sky130_fd_io__tk_em1o
XI38 net144 net134 sky130_fd_io__tk_em1o
XI32 net144 net132 sky130_fd_io__tk_em1o
XI83<1> net106<0> vref_nng sky130_fd_io__tk_em1o
XI83<0> net106<1> vref_nng sky130_fd_io__tk_em1o
XI82 net129 net128 sky130_fd_io__tk_em1o
XI98 net142 net126 sky130_fd_io__tk_em1o
XI30 net144 vgnd_io sky130_fd_io__tk_tie_r_out_esd
XI104 net142 vgnd_io sky130_fd_io__tk_tie_r_out_esd
XI81 net245 net152 sky130_fd_io__sio_pudrvr_esd_res
XI79 net151 net160 sky130_fd_io__sio_pudrvr_esd_res
XI80 net128 net148 sky130_fd_io__sio_pudrvr_esd_res
XI78 net128 net146 sky130_fd_io__sio_pudrvr_esd_res
Xresd net110 net162 sky130_fd_io__res250only_small
Xpsw pu_h_n<1> pghs_h pug<1> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<6> net148 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<5> net148 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<4> net148 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<3> net148 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<2> net146 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<1> net146 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<0> net146 pug<1> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<9> net162 pug<0> net196 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI73 pu_h_n<0> pghs_h pug<0> vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP2<2> net122 net184 vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<8> net160 pug<0> net184 vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpdrvr0<7> net152 pug<0> vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=20.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP2<0> net184 net184 vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP2<1> net196 net184 vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMP2<3> net140 net184 vcc_io vpb_drvr sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<13> net221 net138 pad vgnd_io sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<14> net221 net126 pad vgnd_io sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnsw pug<1> nghs_h pu_h_n<1> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<9> net253<0> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<8> net253<1> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<7> net253<2> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<6> net253<3> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<5> net253<4> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<2> net249 net134 pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<4> net245 vref_int net244 pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<3> net249 net112 pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI74 pug<0> nghs_h pu_h_n<0> vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI54<4> net244 drvhi_h pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI54<5> net244 drvhi_h pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<1> net129 net106<0> pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM<0> net129 net106<1> pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<13> net225<0> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<12> net225<1> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<11> net225<2> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XMa<10> net225<3> net132 pad pad sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__sio_pudrvr_reg drvhi_h en_hicc fb_in fb_out nghs_h pad pghs_h 
+ pu_h_n<1> pu_h_n<0> puen_reg_h pug<1> pug<0> refleak_bias slow_h_n vcc_io 
+ vgnd vgnd_io voutref vpb_drvr vpwr_ka vreg_en_h
*.PININFO drvhi_h:I en_hicc:I fb_in:I nghs_h:I pghs_h:I pu_h_n<1>:I 
*.PININFO pu_h_n<0>:I puen_reg_h:I refleak_bias:I slow_h_n:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I voutref:I vpb_drvr:I vpwr_ka:I vreg_en_h:I fb_out:O pad:B 
*.PININFO pug<1>:B pug<0>:B
XI425 net78 net87 net89 net79 vgnd vpwr_ka vpwr_ka 
+ sky130_fd_io__sio_in_ctl_ls_out_reg
XI429 vreg_en_h net87 sky130_fd_io__tk_em1o_b
XI430 puen_reg_h net87 sky130_fd_io__tk_em1s
Xleak_bias nbias vgnd vpwr_ka vpwr_ka net89 sky130_fd_io__sio_opamp_biasgen_reg
Xreg_opamp en_hicc fb_in fb_out refleak_bias vcc_io vgnd voutref net87 net78 
+ sky130_fd_io__sio_pudrvr_reg_opamp_c
Xleak_inst pad pu_h_n<1> nbias vcc_io vgnd sky130_fd_io__sio_pudrvr_reg_leak
Xcsw_inst drvhi_h puen_reg_h slow_h_n vcc_io vgnd vpwr_ka vref_nng fb_out 
+ sky130_fd_io__sio_pudrvr_reg_csw
Xpu_inst drvhi_h nghs_h pad pghs_h pu_h_n<1> pu_h_n<0> pug<1> pug<0> vcc_io 
+ vgnd vgnd_io vpb_drvr fb_out vref_nng sky130_fd_io__sio_pudrvr_reg_pu
.ENDS

.SUBCKT sky130_fd_io__sio_odrvr_sub drvhi_h od_h oe_hs_h pad pd_h<4> pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pu_h_n<5> pu_h_n<4> pu_h_n<3> pu_h_n<2> pu_h_n<1> 
+ pu_h_n<0> puen_reg_h refleak_bias slow_h_n tie_lo_esd vcc_io vgnd vgnd_io 
+ voutref vpwr_ka vreg_en_h
*.PININFO drvhi_h:I od_h:I oe_hs_h:I pd_h<4>:I pd_h<3>:I pd_h<2>:I pd_h<1>:I 
*.PININFO pd_h<0>:I pu_h_n<5>:I pu_h_n<4>:I pu_h_n<3>:I pu_h_n<2>:I 
*.PININFO pu_h_n<1>:I pu_h_n<0>:I puen_reg_h:I refleak_bias:I slow_h_n:I 
*.PININFO vcc_io:I vgnd:I vgnd_io:I voutref:I vpwr_ka:I vreg_en_h:I pad:O 
*.PININFO tie_lo_esd:O
XI122<4> pd_h<4> pghs_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI122<3> pd_h<3> pghs_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI122<2> pd_h<2> pghs_h vgnd_io vgnd_io sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=20.0 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xhotswap tie_lo_esd od_h oe_hs_h p2g pad pghs_h pug_h<5> pug_h<4> pug_h<3> 
+ pug_h<2> pug_h<1> pug_h<0> vcc_io vcc_io_soft vgnd vpb_drvr vcc_io 
+ sky130_fd_io__sio_hotswap
Xrtie_hi vcc_io tie_hi sky130_fd_io__sio_tk_tie_r
Xodrvr tie_hi p2g pad pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<3> pug_h<2> pug_h<1> pug_h<0> tie_lo_esd 
+ vcc_io vcc_io_soft vgnd vgnd_io vpb_drvr sky130_fd_io__sio_odrvr_nonreg
Xpudrvr_reg drvhi_h vcc_io_soft vref_int vref_int tie_hi pad pghs_h pu_h_n<5> 
+ pu_h_n<4> puen_reg_h pug_h<5> pug_h<4> refleak_bias slow_h_n vcc_io vgnd 
+ vgnd_io voutref vpb_drvr vpwr_ka vreg_en_h sky130_fd_io__sio_pudrvr_reg
.ENDS

.SUBCKT sky130_fd_io__sio_odrvr drvhi_h od_h oe_hs_h pad pd_h<4> pd_h<3> pd_h<2> 
+ pd_h<1> pd_h<0> pu_h_n<5> pu_h_n<4> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> 
+ puen_reg_h refleak_bias slow_h_n tie_lo_esd vcc_io vgnd vgnd_io voutref 
+ vpwr_ka vreg_en_h
*.PININFO drvhi_h:I od_h:I oe_hs_h:I pd_h<4>:I pd_h<3>:I pd_h<2>:I pd_h<1>:I 
*.PININFO pd_h<0>:I pu_h_n<5>:I pu_h_n<4>:I pu_h_n<3>:I pu_h_n<2>:I 
*.PININFO pu_h_n<1>:I pu_h_n<0>:I puen_reg_h:I refleak_bias:I slow_h_n:I 
*.PININFO vcc_io:I vgnd:I vgnd_io:I voutref:I vpwr_ka:I vreg_en_h:I pad:O 
*.PININFO tie_lo_esd:O
Xbondpad pad vgnd_io sky130_fd_io__com_pad
Xodrv_sub drvhi_h od_h oe_hs_h pad pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pu_h_n<5> pu_h_n<4> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_reg_h 
+ refleak_bias slow_h_n tie_lo_esd vcc_io vgnd vgnd_io voutref vpwr_ka 
+ vreg_en_h sky130_fd_io__sio_odrvr_sub
.ENDS

.SUBCKT sky130_fd_io__sio_opath din dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hld_i_ovr_h hld_i_vpwr od_h oe_n pad refleak_bias slow 
+ tie_lo_esd vcc_io vgnd vgnd_io voutref vpwr vpwr_ka vreg_en
*.PININFO din:I dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I 
*.PININFO dm_h_n<0>:I hld_i_h_n:I hld_i_ovr_h:I hld_i_vpwr:I od_h:I oe_n:I 
*.PININFO refleak_bias:I slow:I vcc_io:I vgnd:I vgnd_io:I voutref:I vpwr:I 
*.PININFO vpwr_ka:I vreg_en:I pad:O tie_lo_esd:O
Xopath din dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h 
+ hld_i_h_n hld_i_ovr_h hld_i_vpwr od_h oe_hs_h oe_n pd_h<4> pd_h<3> pd_h<2> 
+ pd_h<1> pd_h<0> pu_h_n<5> pu_h_n<4> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> 
+ puen_reg_h slow slow_h_n vcc_io vgnd vgnd_io vpwr vpwr_ka vreg_en vreg_en_h 
+ sky130_fd_io__sio_opath_sub
Xodrvr drvhi_h od_h oe_hs_h pad pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pu_h_n<5> pu_h_n<4> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_reg_h 
+ refleak_bias slow_h_n tie_lo_esd vcc_io vgnd vgnd_io voutref vpwr_ka 
+ vreg_en_h sky130_fd_io__sio_odrvr
.ENDS

.SUBCKT sky130_fd_io__top_sio dm<2> dm<1> dm<0> enable_h hld_h_n hld_ovr ibuf_sel 
+ in in_h inp_dis oe_n out pad pad_a_esd_0_h pad_a_esd_1_h pad_a_noesd_h 
+ refleak_bias slow tie_lo_esd vccd vcchib vddio vddio_q vinref voutref 
+ vreg_en vssd vssio vssio_q vtrip_sel
*.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I hld_h_n:I hld_ovr:I ibuf_sel:I 
*.PININFO inp_dis:I oe_n:I out:I refleak_bias:I slow:I vinref:I voutref:I 
*.PININFO vreg_en:I vtrip_sel:I in:O in_h:O tie_lo_esd:O pad:B pad_a_esd_0_h:B 
*.PININFO pad_a_esd_1_h:B pad_a_noesd_h:B vccd:B vcchib:B vddio:B vddio_q:B 
*.PININFO vssd:B vssio:B vssio_q:B
Xipath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> ibuf_sel_h 
+ ibuf_sel_h_n inp_dis_h inp_dis_h_n in in_h pad tie_lo_esd vddio vddio_q vssd 
+ vinref vcchib vcchib trip_sel_h trip_sel_h_n sky130_fd_io__sio_ipath_tsg4
Xcom_ctl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> enable_h hld_h_n hld_i_h_n hld_i_ovr_h hld_i_vpwr hld_ovr ibuf_sel 
+ ibuf_sel_h ibuf_sel_h_n inp_dis inp_dis_h inp_dis_h_n net94 vddio_q vssd 
+ vccd vtrip_sel trip_sel_h trip_sel_h_n sky130_fd_io__sio_ctl
XI70 pad_a_esd_0_h pad sky130_fd_io__sio_res250only_small_esd
XI103 pad_a_esd_1_h pad sky130_fd_io__sio_res250only_small_esd
Xopath out dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_ovr_h hld_i_vpwr net94 oe_n pad refleak_bias slow tie_lo_esd vddio 
+ vssd vssio voutref vccd vcchib vreg_en sky130_fd_io__sio_opath
RI71 pad pad_a_noesd_h sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__top_sio_macro amuxbus_a amuxbus_b dft_refgen dm0<2> dm0<1> 
+ dm0<0> dm1<2> dm1<1> dm1<0> enable_h enable_vdda_h hld_h_n<1> hld_h_n<0> 
+ hld_h_n_refgen hld_ovr<1> hld_ovr<0> ibuf_sel<1> ibuf_sel<0> ibuf_sel_refgen 
+ in<1> in<0> in_h<1> in_h<0> inp_dis<1> inp_dis<0> oe_n<1> oe_n<0> out<1> 
+ out<0> pad<1> pad<0> pad_a_esd_0_h<1> pad_a_esd_0_h<0> pad_a_esd_1_h<1> 
+ pad_a_esd_1_h<0> pad_a_noesd_h<1> pad_a_noesd_h<0> slow<1> slow<0> 
+ tie_lo_esd<1> tie_lo_esd<0> vccd vcchib vdda vddio vddio_q vinref_dft 
+ voh_sel<2> voh_sel<1> voh_sel<0> vohref voutref_dft vref_sel<1> vref_sel<0> 
+ vreg_en<1> vreg_en<0> vreg_en_refgen vssa vssd vssio vssio_q vswitch 
+ vtrip_sel<1> vtrip_sel<0> vtrip_sel_refgen
*.PININFO dft_refgen:I dm0<2>:I dm0<1>:I dm0<0>:I dm1<2>:I dm1<1>:I dm1<0>:I 
*.PININFO enable_h:I enable_vdda_h:I hld_h_n<1>:I hld_h_n<0>:I 
*.PININFO hld_h_n_refgen:I hld_ovr<1>:I hld_ovr<0>:I ibuf_sel<1>:I 
*.PININFO ibuf_sel<0>:I ibuf_sel_refgen:I inp_dis<1>:I inp_dis<0>:I oe_n<1>:I 
*.PININFO oe_n<0>:I out<1>:I out<0>:I slow<1>:I slow<0>:I voh_sel<2>:I 
*.PININFO voh_sel<1>:I voh_sel<0>:I vohref:I vref_sel<1>:I vref_sel<0>:I 
*.PININFO vreg_en<1>:I vreg_en<0>:I vreg_en_refgen:I vtrip_sel<1>:I 
*.PININFO vtrip_sel<0>:I vtrip_sel_refgen:I in<1>:O in<0>:O in_h<1>:O 
*.PININFO in_h<0>:O tie_lo_esd<1>:O tie_lo_esd<0>:O amuxbus_a:B amuxbus_b:B 
*.PININFO pad<1>:B pad<0>:B pad_a_esd_0_h<1>:B pad_a_esd_0_h<0>:B 
*.PININFO pad_a_esd_1_h<1>:B pad_a_esd_1_h<0>:B pad_a_noesd_h<1>:B 
*.PININFO pad_a_noesd_h<0>:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B 
*.PININFO vinref_dft:B voutref_dft:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
XREFGEN amuxbus_a amuxbus_b dft_refgen enable_h enable_vdda_h hld_h_n_refgen 
+ ibuf_sel_refgen refleak_bias vccd vcchib vdda vddio vddio_q vinref 
+ vinref_dft voh_sel<2> voh_sel<1> voh_sel<0> vohref voutref voutref_dft 
+ vref_sel<1> vref_sel<0> vreg_en_refgen vssa vssd vssio vssio_q vswitch 
+ vtrip_sel_refgen sky130_fd_io__top_refgen_new
XSIO_PAIR<1> dm1<2> dm1<1> dm1<0> enable_h hld_h_n<1> hld_ovr<1> ibuf_sel<1> 
+ in<1> in_h<1> inp_dis<1> oe_n<1> out<1> pad<1> pad_a_esd_0_h<1> 
+ pad_a_esd_1_h<1> pad_a_noesd_h<1> refleak_bias slow<1> tie_lo_esd<1> vccd 
+ vcchib vddio vddio_q vinref voutref vreg_en<1> vssd vssio vssio_q 
+ vtrip_sel<1> sky130_fd_io__top_sio
XSIO_PAIR<0> dm0<2> dm0<1> dm0<0> enable_h hld_h_n<0> hld_ovr<0> ibuf_sel<0> 
+ in<0> in_h<0> inp_dis<0> oe_n<0> out<0> pad<0> pad_a_esd_0_h<0> 
+ pad_a_esd_1_h<0> pad_a_noesd_h<0> refleak_bias slow<0> tie_lo_esd<0> vccd 
+ vcchib vddio vddio_q vinref voutref vreg_en<0> vssd vssio vssio_q 
+ vtrip_sel<0> sky130_fd_io__top_sio
.ENDS

.SUBCKT sky130_fd_io__tp1_res a b
*.PININFO a:B b:B
XRI21 a net27 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI0 net27 net23 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI1 net25 net17 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI2 net23 net25 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI3 net21 net19 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI4 net19 b sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI5 net17 net15 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI10 net15 net13 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
XRI9 net13 net21 sky130_fd_pr__res_generic_po m=1 w=0.4 l=112
.ENDS

.SUBCKT sky130_fd_io__tp1_div en_tp1 force_tp1 tp1 tp1_div vnb vssd
*.PININFO en_tp1:I force_tp1:I tp1:I vnb:I vssd:I tp1_div:O
XRESHI<6> tp1 tp1_res<5> sky130_fd_io__tp1_res
XRESHI<5> tp1_res<5> tp1_res<4> sky130_fd_io__tp1_res
XRESHI<4> tp1_res<4> tp1_res<3> sky130_fd_io__tp1_res
XRESHI<3> tp1_res<3> tp1_res<2> sky130_fd_io__tp1_res
XRESHI<2> tp1_res<2> tp1_res<1> sky130_fd_io__tp1_res
XRESHI<1> tp1_res<1> tp1_div_int sky130_fd_io__tp1_res
XRESLO tp1_div_int tp1_sw sky130_fd_io__tp1_res
XM0 tp1_sw en_tp1 vssd vnb sky130_fd_pr__nfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 sa=2 sb=2.5 sd=0.28 
+ topography=normal area=0.063 perim=1.14
XM2 tp1_div_int en_tp1 tp1_div vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=2 sb=2.5 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XM1 tp1_div_int force_tp1 vssd vnb sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=2 sb=2.5 
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__res250only pad rout
*.PININFO pad:B rout:B
XRI175 net12 net16 sky130_fd_pr__res_generic_po m=1 w=4 l=20.195
XRI229 net16 rout sky130_fd_pr__res_generic_po m=1 w=4 l=0.17
XRI228 pad net12 sky130_fd_pr__res_generic_po m=1 w=4 l=0.17
RI237<1> net16 rout sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI237<2> net16 rout sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI234<1> pad net12 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
RI234<2> pad net12 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__signal_40_sym_hv_2k_dnwl_aup1_b body g<5> g<4> g<3> g<2> g<1> 
+ g<0> gate<9> gate<8> gate<7> gate<6> gate<5> gate<4> gate<3> gate<2> gate<1> 
+ gate<0> nwellRing pad<4> pad<3> pad<2> pad<1> pad<0>
*.PININFO gate<9>:I gate<8>:I gate<7>:I gate<6>:I gate<5>:I gate<4>:I 
*.PININFO gate<3>:I gate<2>:I gate<1>:I gate<0>:I nwellRing:I body:B g<5>:B 
*.PININFO g<4>:B g<3>:B g<2>:B g<1>:B g<0>:B pad<4>:B pad<3>:B pad<2>:B 
*.PININFO pad<1>:B pad<0>:B
XesdNfet4<1> pad<4> gate<9> g<5> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet4<0> pad<4> gate<8> g<4> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet2<1> pad<2> gate<5> g<3> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet2<0> pad<2> gate<4> g<2> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet3<1> pad<3> gate<7> g<4> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet3<0> pad<3> gate<6> g<3> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet1<1> pad<1> gate<3> g<2> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet1<0> pad<1> gate<2> g<1> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet0<1> pad<0> gate<1> g<1> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XesdNfet0<0> pad<0> gate<0> g<0> body sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
RI8 nwellRing net59 sky130_fd_pr__res_generic_m1 l=0.01 w=0.5
.ENDS

.SUBCKT sky130_fd_io__top_tp1 amuxbus_a amuxbus_b en_tp1 tp1 tp1_div tp1_out vccd 
+ vcchib vdda vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO en_tp1:I tp1_div:O amuxbus_a:B amuxbus_b:B tp1:B tp1_out:B vccd:B 
*.PININFO vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B 
*.PININFO vswitch:B
XTP1_DIV en_tp1 vssd tp1_out tp1_div vssd vssd sky130_fd_io__tp1_div
XRESD tp1 tp1_out sky130_fd_io__res250only
XESD vssio vssio vssio vssio vssio vssio vssio net68 net68 net68 net68 net68 
+ net68 net68 net68 net68 net68 vddio tp1 tp1 tp1 tp1 tp1 
+ sky130_fd_io__signal_40_sym_hv_2k_dnwl_aup1_b
XRR1 vssio net68 sky130_fd_pr__res_generic_po m=1 w=0.5 l=10.2
.ENDS

.SUBCKT sky130_fd_io__tp2_res a b
*.PININFO a:B b:B
XRR1<8> a n<7> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<7> n<7> n<6> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<6> n<6> n<5> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<5> n<5> n<4> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<4> n<4> n<3> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<3> n<3> n<2> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<2> n<2> n<1> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<1> n<1> n<0> sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
XRR1<0> n<0> b sky130_fd_pr__res_generic_po m=1 w=0.4 l=87
.ENDS

.SUBCKT sky130_fd_io__tp2_ls in out vgnd vhv
*.PININFO in:I vgnd:I vhv:I out:O
XM5 outb out vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM1 ainv in vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XM4 out outb vhv vhv sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM0 ainv in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM2 out ainv vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM3 outb in vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__tp2_inv_1 A Y vgnd vnb vpb vpwr
*.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XMIP1 Y A vpwr vpb sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
XMIN1 Y A vgnd vnb sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__tp2_div en_tp2 force_tp2 tp2 tp2_div vccd vio vssd
*.PININFO en_tp2:I force_tp2:I tp2:I vccd:I vio:I vssd:I tp2_div:O
XRESHI rtop tp2div sky130_fd_io__tp2_res
XRESLO<8> tp2 tp2_res<7> sky130_fd_io__tp2_res
XRESLO<7> tp2_res<7> tp2_res<6> sky130_fd_io__tp2_res
XRESLO<6> tp2_res<6> tp2_res<5> sky130_fd_io__tp2_res
XRESLO<5> tp2_res<5> tp2_res<4> sky130_fd_io__tp2_res
XRESLO<4> tp2_res<4> tp2_res<3> sky130_fd_io__tp2_res
XRESLO<3> tp2_res<3> tp2_res<2> sky130_fd_io__tp2_res
XRESLO<2> tp2_res<2> tp2_res<1> sky130_fd_io__tp2_res
XRESLO<1> tp2_res<1> tp2_div_int sky130_fd_io__tp2_res
XLEVSHIFT en_tp2 en_tp2_hv vssd vio sky130_fd_io__tp2_ls
XU1 force_tp2 forceb_tp2 vssd vssd vccd vccd sky130_fd_io__tp2_inv_1
XU2 en_tp2 enb_tp2 vssd vssd vccd vccd sky130_fd_io__tp2_inv_1
XU3 enb_tp2 en_tp2_buf vssd vssd vccd vccd sky130_fd_io__tp2_inv_1
XM2 tp2_div en_tp2_hv pullup vssd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM3 pullup enb_tp2 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM0 tp2div en_tp2_buf tp2_div_int tp2div sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM6 en_tp2_hv enb_tp2 vssd vssd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM1 tp2div enb_tp2 pullup pullup sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XM4 rtop enb_tp2 vccd vccd sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XM5 rtop forceb_tp2 vccd vccd sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__top_tp2 amuxbus_a amuxbus_b en_tp2 tp2 tp2_div tp2_out vccd 
+ vcchib vdda vddio vddio_q vneg vssa vssd vssio vssio_q vswitch
*.PININFO en_tp2:I tp2_div:O amuxbus_a:B amuxbus_b:B tp2:B tp2_out:B vccd:B 
*.PININFO vcchib:B vdda:B vddio:B vddio_q:B vneg:B vssa:B vssd:B vssio:B 
*.PININFO vssio_q:B vswitch:B
XTP2_DIV en_tp2 vssd tp2_out tp2_div vccd vddio vssd sky130_fd_io__tp2_div
XESD vneg vssio vssio vssio vssio vssio vssio net73 net73 net73 net73 net73 
+ net73 net73 net73 net73 net73 vddio tp2 tp2 tp2 tp2 tp2 
+ sky130_fd_io__signal_40_sym_hv_2k_dnwl_aup1_b
XRI18 vneg net73 sky130_fd_pr__res_generic_po m=1 w=0.5 l=10.2
XRESD tp2 tp2_out sky130_fd_io__res250only
.ENDS

.SUBCKT sky130_fd_io__top_tp3 tp3 tp3_out vddd vssd
*.PININFO tp3:B tp3_out:B vddd:B vssd:B
XRESD tp3 tp3_out sky130_fd_io__res250only
XESD vssd vssd vssd vssd vssd vssd vssd net22 net22 net22 net22 net22 net22 
+ net22 net22 net22 net22 vddd tp3 tp3 tp3 tp3 tp3 
+ sky130_fd_io__signal_40_sym_hv_2k_dnwl_aup1_b
XRR1 vssd net22 sky130_fd_pr__res_generic_po m=1 w=0.5 l=10.2
.ENDS

.SUBCKT sky130_fd_io__xres_ipath in_h in_vt out out_h vcchib vddio_q vssd
*.PININFO in_h:I in_vt:I out:O out_h:O vcchib:B vddio_q:B vssd:B
Xgpio_inbuf vddio_q in_h in_vt out_gpio_h net40 vddio_q vssd vcchib vddio_q 
+ sky130_fd_io__gpio_in_buf
Xrcfilt out_gpio_h out_rcfilt_h vddio_q vssd sky130_fd_io__xres_rcfilter_lpf
Xhyst_buf out_rcfilt_h out_hysbuf_h vddio_q vssd sky130_fd_io__xres_inv_hys
Xhv_lv_ls out_hysbuf_h net56 out vcchib vddio_q vssd sky130_fd_io__xres_hvlv_ls
Xhv_drv1 out_hysbuf_h out_h_n vssd vddio_q sky130_fd_io__hvsbt_inv_x1
Xhv_drv2 out_h_n out_h vssd vddio_q sky130_fd_io__hvsbt_inv_x4
.ENDS

.SUBCKT sky130_fd_io__top_xres_2 amuxbus_a amuxbus_b out out_h pad vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO out:O out_h:O amuxbus_a:B amuxbus_b:B pad:B vccd:B vcchib:B vdda:B 
*.PININFO vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xweakpullup pad vddio vssd sky130_fd_io__xres_wpu
Xxresesd in_h in_vt pad vddio vssd vssio sky130_fd_io__xres_esd
Xibuf in_h in_vt out out_h vcchib vddio_q vssd sky130_fd_io__xres_ipath
.ENDS

.SUBCKT sky130_fd_io__gpio_in_buf_xres2v2 in_h in_vt out_h out_h_n vcc_io vgnd vpwr
*.PININFO in_h:I in_vt:I vcc_io:I vgnd:I vpwr:I out_h:O out_h_n:O
XI49 vcc_io tie_hi_esd sky130_fd_io__tk_tie_r_out_esd
XI599 vpwr net056 sky130_fd_io__tk_tie_r_out_esd
XI596 out_a net115 sky130_fd_io__tk_em1s
Xttl_pd_op net077 net118 sky130_fd_io__tk_em1o
XI576 tie_hi_esd vtrip_sel_h vgnd vcc_io sky130_fd_io__hvsbt_inv_x1
Xpd2 net134 out_a vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1_mid_nat net130 net056 net103 vgnd sky130_fd_pr__nfet_05v0_nvt m=4 w=1.00 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpd_hrng net118 in_vt net117 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=3.00 l=1.00 mult=1 sa=0.265 
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpden_1 net117 tie_hi_esd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=12 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpd1 net118 in_h net117 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI585 net115 net115 out_a vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI574 net118 out_a net137 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI598 net118 out_a vcc_io vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI592 out_h out_h_n vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI584 net103 net103 net115 vgnd sky130_fd_pr__nfet_05v0_nvt m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI571 net118 out_a vcc_io vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI597 net118 out_a net137 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI570 out_a in_h net118 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI595 net077 in_vt net117 vgnd sky130_fd_pr__nfet_g5v0d10v5 m=8 w=3.00 l=1.00 mult=1 sa=0.265 sb=0.265 
+ sd=0.28 topography=normal area=0.063 perim=1.14
XI589 out_h_n net134 vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xdis_trip_sel1 in_vt tie_hi_esd vgnd vgnd sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu2 net134 out_a vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1 net169 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpuen_2 out_a tie_hi_esd vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu1_midopt net169 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI567 net130 in_h net169 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI568 vgnd out_a net169 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI590 out_h_n net134 vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI579 net153 in_h vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI578 out_a in_h net153 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI593 out_h out_h_n vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI577 out_a vtrip_sel_h net130 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI582 vgnd out_a net153 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI575 vcc_io vtrip_sel_h net137 vcc_io sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS

.SUBCKT sky130_fd_io__xres_ipath_xres2v2 in_h in_vt out out_h vcchib vddio_q vssd
*.PININFO in_h:I in_vt:I out:O out_h:O vcchib:B vddio_q:B vssd:B
XI35 out net018 vssd vssd sky130_fd_pr__nfet_01v8 m=8 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI34 net018 net061 vssd vssd sky130_fd_pr__nfet_01v8 m=2 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI32 net018 net061 vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI33 out net018 vcchib vcchib sky130_fd_pr__pfet_01v8_hvt m=4 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xgpio_inbuf in_h in_vt out_gpio_h net40 vddio_q vssd vcchib 
+ sky130_fd_io__gpio_in_buf_xres2v2
Xrcfilt out_gpio_h out_rcfilt_h vddio_q vssd sky130_fd_io__xres_rcfilter_lpf
Xhyst_buf out_rcfilt_h out_hysbuf_h vddio_q vssd sky130_fd_io__xres_inv_hys
Xhv_lv_ls out_hysbuf_h net56 net061 vcchib vddio_q vssd sky130_fd_io__xres_hvlv_ls
Xhv_drv1 out_hysbuf_h out_h_n vssd vddio_q sky130_fd_io__hvsbt_inv_x1
Xhv_drv2 out_h_n out_h vssd vddio_q sky130_fd_io__hvsbt_inv_x4
.ENDS

.SUBCKT sky130_fd_io__top_xres2v2 amuxbus_a amuxbus_b pad vccd vcchib vdda vddio 
+ vddio_q vssa vssd vssio vssio_q vswitch xres_h_n xres_n
*.PININFO xres_h_n:O xres_n:O amuxbus_a:B amuxbus_b:B pad:B vccd:B vcchib:B 
*.PININFO vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xesd_res pad net35 sky130_fd_io__res250only_small
Xxresesd in_h in_vt pad vddio vssd vssio sky130_fd_io__xres_esd
Xweakpullup net35 vddio vssd sky130_fd_io__xres_wpu
Xibuf in_h in_vt xres_n xres_h_n vcchib vddio_q vssd 
+ sky130_fd_io__xres_ipath_xres2v2
.ENDS

.SUBCKT sky130_fd_io__top_xres3v2 amuxbus_a amuxbus_b pad pad_a_esd_h tie_weak_hi_h 
+ vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q vswitch xres_h_n 
+ xres_n
*.PININFO xres_h_n:O xres_n:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_h:B 
*.PININFO tie_weak_hi_h:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B 
*.PININFO vssd:B vssio:B vssio_q:B vswitch:B
Xesd_res pad pad_a_esd_h sky130_fd_io__res250only_small
Xibuf in_h in_vt xres_n xres_h_n vcchib vddio_q vssd 
+ sky130_fd_io__xres_ipath_xres2v2
Xweakpullup tie_weak_hi_h vddio vssd sky130_fd_io__xres_wpu
Xxresesd in_h in_vt pad vddio vssd vssio sky130_fd_io__xres_esd
.ENDS

.SUBCKT sky130_fd_io__top_xres amuxbus_a amuxbus_b out out_h pad vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO out:O out_h:O amuxbus_a:B amuxbus_b:B pad:B vccd:B vcchib:B vdda:B 
*.PININFO vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xweakpullup pad vddio vssd sky130_fd_io__xres_wpu
Xxresesd in_h in_vt pad vddio vssd vssio sky130_fd_io__xres_esd
Xibuf in_h in_vt out out_h vcchib vddio_q vssd sky130_fd_io__xres_ipath
.ENDS
